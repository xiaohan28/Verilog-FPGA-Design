`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/18/2024 05:51:42 PM
// Design Name: 
// Module Name: frame_data
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module start_screen(input frame_rate, input [12:0] pixel_index, output reg [15:0] oled_data);
    reg [15:0] frame_count = 1;
    parameter picture_total_count = 1;
    
    always @ (posedge frame_rate) begin
        frame_count <= (frame_count == picture_total_count - 1) ? 0 : frame_count + 1;
    end
   
    always @ (*) begin
   case (pixel_index)
    0, 1, 2, 3, 4, 5, 6, 7, 8, 9: oled_data = 16'b1111111111111111;
    10, 11, 12, 13, 14, 15, 16, 17, 18, 19: oled_data = 16'b1111111111111111;
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29: oled_data = 16'b1111111111111111;
    30, 31, 32, 33, 34, 35, 36, 37, 38, 39: oled_data = 16'b1111111111111111;
    40, 41, 42, 43, 44, 45, 46, 47, 48, 49: oled_data = 16'b1111111111111111;
    50, 51, 52, 53, 54, 55, 56, 57, 58, 59: oled_data = 16'b1111111111111111;
    60, 61, 62, 63, 64, 65, 66, 67, 68, 69: oled_data = 16'b1111111111111111;
    70, 71, 72, 73, 74, 75, 76, 77, 78, 79: oled_data = 16'b1111111111111111;
    80, 81, 82, 83, 84, 85, 86, 87, 88, 89: oled_data = 16'b1111111111111111;
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99: oled_data = 16'b1111111111111111;
    100, 101, 102, 103, 104, 105, 106, 107, 108, 109: oled_data = 16'b1111111111111111;
    110, 111, 112, 113, 114, 115, 116, 117, 118, 119: oled_data = 16'b1111111111111111;
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129: oled_data = 16'b1111111111111111;
    130, 131, 132, 133, 134, 135, 136, 137, 138, 139: oled_data = 16'b1111111111111111;
    140, 141, 142, 143, 144, 145, 146, 147, 148, 149: oled_data = 16'b1111111111111111;
    150, 151, 152, 153, 154, 155, 156, 157, 158, 159: oled_data = 16'b1111111111111111;
    160, 161, 162, 163, 164, 165, 166, 167, 168, 169: oled_data = 16'b1111111111111111;
    170, 171, 172, 173, 174, 175, 176, 177, 178, 179: oled_data = 16'b1111111111111111;
    180, 181, 182, 183, 184, 185, 186, 187, 188, 189: oled_data = 16'b1111111111111111;
    190, 191, 192, 193, 194, 195, 196, 197, 198, 199: oled_data = 16'b1111111111111111;
    200, 201, 203, 204, 205, 206, 207, 208, 209, 210: oled_data = 16'b1111111111111111;
    213, 214, 215, 216, 217, 219, 220, 221, 222, 223: oled_data = 16'b1111111111111111;
    224, 225, 227, 228, 229, 230, 231, 232, 233, 234: oled_data = 16'b1111111111111111;
    236, 237, 238, 239, 240, 242, 243, 244, 245, 246: oled_data = 16'b1111111111111111;
    247, 248, 249, 250, 251, 252, 253, 254, 255, 256: oled_data = 16'b1111111111111111;
    257, 260, 261, 262, 263, 264, 266, 267, 268, 269: oled_data = 16'b1111111111111111;
    270, 271, 272, 273, 274, 275, 277, 278, 279, 280: oled_data = 16'b1111111111111111;
    281, 282, 283, 284, 285, 286, 287, 288, 289, 290: oled_data = 16'b1111111111111111;
    291, 292, 293, 294, 295, 296, 297, 298, 299, 300: oled_data = 16'b1111111111111111;
    301, 302, 303, 304, 305, 306, 307, 308, 309, 310: oled_data = 16'b1111111111111111;
    311, 312, 313, 314, 315, 316, 317, 318, 319, 320: oled_data = 16'b1111111111111111;
    321, 322, 323, 324, 325, 326, 327, 328, 329, 330: oled_data = 16'b1111111111111111;
    331, 332, 333, 334, 335, 336, 337, 338, 339, 340: oled_data = 16'b1111111111111111;
    341, 342, 343, 344, 345, 346, 347, 348, 349, 350: oled_data = 16'b1111111111111111;
    351, 352, 353, 354, 355, 356, 357, 358, 359, 360: oled_data = 16'b1111111111111111;
    361, 362, 363, 364, 365, 366, 367, 368, 369, 370: oled_data = 16'b1111111111111111;
    371, 372, 373, 374, 375, 376, 377, 378, 379, 380: oled_data = 16'b1111111111111111;
    381, 382, 383, 384, 385, 386, 387, 388, 389, 390: oled_data = 16'b1111111111111111;
    391, 398, 399, 400, 406, 407, 411, 419, 423, 424: oled_data = 16'b1111111111111111;
    425, 429, 430, 436, 441, 442, 447, 453, 454, 458: oled_data = 16'b1111111111111111;
    459, 460, 464, 465, 471, 472, 473, 474, 475, 476: oled_data = 16'b1111111111111111;
    477, 478, 479, 480, 481, 482, 483, 484, 485, 486: oled_data = 16'b1111111111111111;
    487, 494, 496, 503, 507, 515, 519, 525, 532, 543: oled_data = 16'b1111111111111111;
    550, 560, 567, 568, 569, 570, 571, 572, 573, 574: oled_data = 16'b1111111111111111;
    575, 576, 577, 578, 579, 580, 581, 582, 583, 611: oled_data = 16'b1111111111111111;
    664, 665, 666, 667, 668, 669, 670, 671, 672, 673: oled_data = 16'b1111111111111111;
    674, 675, 676, 677, 678, 679, 683, 691, 702, 703: oled_data = 16'b1111111111111111;
    707, 721, 738, 756, 760, 761, 762, 763, 764, 765: oled_data = 16'b1111111111111111;
    766, 767, 768, 769, 770, 771, 772, 773, 775, 783: oled_data = 16'b1111111111111111;
    798, 799, 803, 856, 858, 859, 860, 861, 862, 863: oled_data = 16'b1111111111111111;
    864, 865, 866, 867, 868, 869, 871, 879, 894, 895: oled_data = 16'b1111111111111111;
    899, 903, 952, 954, 955, 956, 957, 958, 959, 960: oled_data = 16'b1111111111111111;
    961, 962, 963, 964, 965, 966, 967, 971, 979, 991: oled_data = 16'b1111111111111111;
    995, 999, 1017, 1018, 1026, 1034, 1035, 1036, 1044, 1048: oled_data = 16'b1111111111111111;
    1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059: oled_data = 16'b1111111111111111;
    1060, 1061, 1062, 1063, 1071, 1075, 1091, 1095, 1113, 1114: oled_data = 16'b1111111111111111;
    1122, 1132, 1140, 1144, 1145, 1146, 1147, 1148, 1149, 1150: oled_data = 16'b1111111111111111;
    1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159, 1166: oled_data = 16'b1111111111111111;
    1167, 1171, 1179, 1187, 1191, 1197, 1198, 1204, 1209, 1210: oled_data = 16'b1111111111111111;
    1218, 1226, 1227, 1228, 1236, 1240, 1242, 1243, 1244, 1245: oled_data = 16'b1111111111111111;
    1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253, 1254, 1255: oled_data = 16'b1111111111111111;
    1262, 1263, 1267, 1271, 1275, 1279, 1283, 1287, 1288, 1289: oled_data = 16'b1111111111111111;
    1293, 1299, 1300, 1301, 1305, 1306, 1310, 1314, 1318, 1322: oled_data = 16'b1111111111111111;
    1323, 1324, 1328, 1332, 1336, 1337, 1338, 1339, 1340, 1341: oled_data = 16'b1111111111111111;
    1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351: oled_data = 16'b1111111111111111;
    1352, 1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361: oled_data = 16'b1111111111111111;
    1362, 1363, 1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371: oled_data = 16'b1111111111111111;
    1372, 1373, 1374, 1375, 1376, 1377, 1378, 1379, 1380, 1381: oled_data = 16'b1111111111111111;
    1382, 1383, 1384, 1385, 1386, 1387, 1388, 1389, 1390, 1391: oled_data = 16'b1111111111111111;
    1392, 1393, 1394, 1395, 1396, 1397, 1398, 1399, 1400, 1401: oled_data = 16'b1111111111111111;
    1402, 1403, 1404, 1405, 1406, 1407, 1408, 1409, 1410, 1411: oled_data = 16'b1111111111111111;
    1412, 1413, 1414, 1415, 1416, 1417, 1418, 1419, 1420, 1421: oled_data = 16'b1111111111111111;
    1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429, 1430, 1431: oled_data = 16'b1111111111111111;
    1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440, 1441: oled_data = 16'b1111111111111111;
    1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451: oled_data = 16'b1111111111111111;
    1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461: oled_data = 16'b1111111111111111;
    1462, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471: oled_data = 16'b1111111111111111;
    1472, 1473, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481: oled_data = 16'b1111111111111111;
    1482, 1483, 1484, 1485, 1486, 1487, 1488, 1489, 1490, 1491: oled_data = 16'b1111111111111111;
    1492, 1493, 1494, 1495, 1496, 1497, 1498, 1499, 1500, 1501: oled_data = 16'b1111111111111111;
    1502, 1503, 1504, 1505, 1506, 1507, 1508, 1509, 1510, 1511: oled_data = 16'b1111111111111111;
    1512, 1513, 1514, 1515, 1516, 1517, 1518, 1519, 1520, 1521: oled_data = 16'b1111111111111111;
    1522, 1523, 1524, 1525, 1526, 1527, 1528, 1529, 1530, 1531: oled_data = 16'b1111111111111111;
    1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539, 1540, 1541: oled_data = 16'b1111111111111111;
    1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550, 1551: oled_data = 16'b1111111111111111;
    1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561: oled_data = 16'b1111111111111111;
    1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571: oled_data = 16'b1111111111111111;
    1572, 1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581: oled_data = 16'b1111111111111111;
    1582, 1583, 1584, 1585, 1586, 1587, 1588, 1589, 1590, 1591: oled_data = 16'b1111111111111111;
    1592, 1593, 1594, 1595, 1596, 1597, 1598, 1599, 1600, 1601: oled_data = 16'b1111111111111111;
    1602, 1603, 1604, 1605, 1606, 1607, 1608, 1609, 1610, 1611: oled_data = 16'b1111111111111111;
    1612, 1613, 1614, 1615, 1616, 1617, 1618, 1619, 1620, 1621: oled_data = 16'b1111111111111111;
    1622, 1623, 1624, 1625, 1626, 1627, 1628, 1629, 1630, 1631: oled_data = 16'b1111111111111111;
    1632, 1633, 1634, 1635, 1636, 1637, 1638, 1639, 1640, 1641: oled_data = 16'b1111111111111111;
    1642, 1643, 1644, 1645, 1646, 1647, 1648, 1649, 1650, 1651: oled_data = 16'b1111111111111111;
    1652, 1653, 1654, 1655, 1656, 1657, 1658, 1659, 1660, 1661: oled_data = 16'b1111111111111111;
    1662, 1663, 1664, 1665, 1666, 1667, 1668, 1669, 1670, 1671: oled_data = 16'b1111111111111111;
    1672, 1673, 1674, 1675, 1676, 1677, 1678, 1679, 1680, 1681: oled_data = 16'b1111111111111111;
    1682, 1683, 1684, 1685, 1686, 1687, 1688, 1689, 1690, 1691: oled_data = 16'b1111111111111111;
    1692, 1693, 1694, 1695, 1696, 1697, 1698, 1699, 1700, 1701: oled_data = 16'b1111111111111111;
    1702, 1703, 1704, 1709, 1710, 1711, 1712, 1713, 1720, 1721: oled_data = 16'b1111111111111111;
    1722, 1723, 1724, 1725, 1726, 1727, 1728, 1729, 1730, 1731: oled_data = 16'b1111111111111111;
    1732, 1733, 1734, 1735, 1736, 1737, 1738, 1739, 1740, 1741: oled_data = 16'b1111111111111111;
    1742, 1743, 1744, 1745, 1746, 1747, 1748, 1749, 1750, 1751: oled_data = 16'b1111111111111111;
    1752, 1753, 1754, 1755, 1756, 1757, 1758, 1759, 1760, 1761: oled_data = 16'b1111111111111111;
    1762, 1763, 1764, 1765, 1766, 1767, 1768, 1769, 1770, 1771: oled_data = 16'b1111111111111111;
    1772, 1773, 1774, 1775, 1776, 1777, 1778, 1779, 1780, 1781: oled_data = 16'b1111111111111111;
    1782, 1783, 1784, 1785, 1786, 1787, 1788, 1789, 1790, 1791: oled_data = 16'b1111111111111111;
    1792, 1793, 1794, 1795, 1796, 1797, 1798, 1799, 1806, 1807: oled_data = 16'b1111111111111111;
    1817, 1818, 1819, 1820, 1821, 1822, 1823, 1824, 1825, 1826: oled_data = 16'b1111111111111111;
    1827, 1828, 1829, 1830, 1831, 1832, 1833, 1834, 1835, 1836: oled_data = 16'b1111111111111111;
    1837, 1838, 1839, 1840, 1841, 1842, 1843, 1844, 1845, 1846: oled_data = 16'b1111111111111111;
    1847, 1848, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856: oled_data = 16'b1111111111111111;
    1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1865, 1866: oled_data = 16'b1111111111111111;
    1867, 1868, 1869, 1870, 1871, 1872, 1873, 1874, 1875, 1876: oled_data = 16'b1111111111111111;
    1877, 1878, 1879, 1880, 1881, 1882, 1883, 1884, 1885, 1886: oled_data = 16'b1111111111111111;
    1887, 1888, 1889, 1890, 1891, 1892, 1893, 1894, 1903, 1904: oled_data = 16'b1111111111111111;
    1913, 1915, 1916, 1917, 1918, 1919, 1920, 1921, 1922, 1923: oled_data = 16'b1111111111111111;
    1924, 1925, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933: oled_data = 16'b1111111111111111;
    1934, 1935, 1936, 1937, 1938, 1939, 1940, 1941, 1942, 1943: oled_data = 16'b1111111111111111;
    1944, 1945, 1946, 1947, 1948, 1949, 1950, 1951, 1952, 1953: oled_data = 16'b1111111111111111;
    1954, 1955, 1956, 1957, 1958, 1959, 1960, 1961, 1962, 1963: oled_data = 16'b1111111111111111;
    1964, 1965, 1966, 1967, 1968, 1969, 1970, 1971, 1972, 1973: oled_data = 16'b1111111111111111;
    1974, 1975, 1976, 1977, 1978, 1979, 1980, 1981, 1982, 1983: oled_data = 16'b1111111111111111;
    1984, 1985, 1986, 1987, 1988, 1989, 2010, 2011, 2012, 2013: oled_data = 16'b1111111111111111;
    2014, 2015, 2016, 2017, 2018, 2019, 2020, 2021, 2022, 2023: oled_data = 16'b1111111111111111;
    2024, 2025, 2026, 2027, 2028, 2029, 2030, 2031, 2032, 2033: oled_data = 16'b1111111111111111;
    2034, 2035, 2036, 2037, 2038, 2039, 2040, 2041, 2042, 2043: oled_data = 16'b1111111111111111;
    2044, 2045, 2046, 2047, 2048, 2049, 2050, 2051, 2052, 2053: oled_data = 16'b1111111111111111;
    2054, 2055, 2056, 2057, 2058, 2059, 2060, 2061, 2062, 2063: oled_data = 16'b1111111111111111;
    2064, 2065, 2066, 2067, 2068, 2069, 2070, 2071, 2072, 2073: oled_data = 16'b1111111111111111;
    2074, 2075, 2076, 2077, 2078, 2079, 2080, 2081, 2082, 2083: oled_data = 16'b1111111111111111;
    2084, 2099, 2107, 2108, 2109, 2110, 2111, 2112, 2113, 2114: oled_data = 16'b1111111111111111;
    2115, 2116, 2117, 2118, 2119, 2120, 2121, 2122, 2123, 2124: oled_data = 16'b1111111111111111;
    2125, 2126, 2127, 2128, 2129, 2130, 2131, 2132, 2133, 2134: oled_data = 16'b1111111111111111;
    2135, 2136, 2137, 2138, 2139, 2140, 2141, 2142, 2143, 2144: oled_data = 16'b1111111111111111;
    2145, 2146, 2147, 2148, 2149, 2150, 2151, 2152, 2153, 2154: oled_data = 16'b1111111111111111;
    2155, 2156, 2157, 2158, 2159, 2160, 2161, 2162, 2163, 2164: oled_data = 16'b1111111111111111;
    2165, 2166, 2167, 2168, 2169, 2170, 2171, 2172, 2173, 2174: oled_data = 16'b1111111111111111;
    2175, 2176, 2177, 2178, 2179, 2180, 2203, 2204, 2205, 2206: oled_data = 16'b1111111111111111;
    2207, 2208, 2209, 2210, 2211, 2212, 2213, 2214, 2215, 2216: oled_data = 16'b1111111111111111;
    2217, 2218, 2219, 2220, 2221, 2222, 2223, 2224, 2225, 2226: oled_data = 16'b1111111111111111;
    2227, 2228, 2229, 2230, 2231, 2232, 2233, 2234, 2235, 2236: oled_data = 16'b1111111111111111;
    2237, 2238, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 2246: oled_data = 16'b1111111111111111;
    2247, 2248, 2249, 2250, 2251, 2252, 2253, 2254, 2255, 2256: oled_data = 16'b1111111111111111;
    2257, 2258, 2259, 2260, 2261, 2262, 2263, 2264, 2265, 2266: oled_data = 16'b1111111111111111;
    2267, 2268, 2269, 2270, 2271, 2272, 2273, 2274, 2275, 2276: oled_data = 16'b1111111111111111;
    2299, 2300, 2301, 2302, 2303, 2304, 2305, 2306, 2307, 2308: oled_data = 16'b1111111111111111;
    2309, 2310, 2311, 2312, 2313, 2314, 2315, 2316, 2317, 2318: oled_data = 16'b1111111111111111;
    2319, 2320, 2321, 2322, 2323, 2324, 2325, 2326, 2327, 2328: oled_data = 16'b1111111111111111;
    2329, 2330, 2331, 2332, 2333, 2334, 2335, 2336, 2337, 2338: oled_data = 16'b1111111111111111;
    2339, 2340, 2341, 2342, 2343, 2344, 2345, 2346, 2347, 2348: oled_data = 16'b1111111111111111;
    2349, 2350, 2351, 2352, 2353, 2354, 2355, 2356, 2357, 2358: oled_data = 16'b1111111111111111;
    2359, 2360, 2361, 2362, 2363, 2364, 2365, 2366, 2367, 2368: oled_data = 16'b1111111111111111;
    2369, 2370, 2371, 2372, 2395, 2396, 2397, 2398, 2399, 2400: oled_data = 16'b1111111111111111;
    2401, 2402, 2403, 2404, 2405, 2406, 2407, 2408, 2409, 2410: oled_data = 16'b1111111111111111;
    2411, 2412, 2413, 2414, 2415, 2416, 2417, 2418, 2419, 2420: oled_data = 16'b1111111111111111;
    2421, 2422, 2423, 2424, 2425, 2426, 2427, 2428, 2429, 2430: oled_data = 16'b1111111111111111;
    2431, 2432, 2433, 2434, 2435, 2436, 2437, 2438, 2439, 2440: oled_data = 16'b1111111111111111;
    2441, 2442, 2443, 2444, 2445, 2446, 2447, 2448, 2449, 2450: oled_data = 16'b1111111111111111;
    2451, 2452, 2453, 2454, 2455, 2456, 2457, 2458, 2459, 2460: oled_data = 16'b1111111111111111;
    2461, 2462, 2463, 2464, 2465, 2466, 2467, 2492, 2493, 2494: oled_data = 16'b1111111111111111;
    2495, 2496, 2497, 2498, 2499, 2500, 2501, 2502, 2503, 2504: oled_data = 16'b1111111111111111;
    2505, 2506, 2507, 2508, 2509, 2510, 2511, 2512, 2513, 2514: oled_data = 16'b1111111111111111;
    2515, 2516, 2517, 2518, 2519, 2520, 2521, 2522, 2523, 2524: oled_data = 16'b1111111111111111;
    2525, 2526, 2527, 2528, 2529, 2530, 2531, 2532, 2533, 2534: oled_data = 16'b1111111111111111;
    2535, 2536, 2537, 2538, 2539, 2540, 2541, 2542, 2543, 2544: oled_data = 16'b1111111111111111;
    2545, 2546, 2547, 2548, 2549, 2550, 2551, 2552, 2553, 2554: oled_data = 16'b1111111111111111;
    2555, 2556, 2557, 2558, 2559, 2560, 2561, 2562, 2563, 2589: oled_data = 16'b1111111111111111;
    2590, 2591, 2592, 2593, 2594, 2595, 2596, 2597, 2598, 2599: oled_data = 16'b1111111111111111;
    2600, 2601, 2602, 2603, 2604, 2605, 2606, 2607, 2608, 2609: oled_data = 16'b1111111111111111;
    2610, 2611, 2612, 2613, 2614, 2615, 2616, 2617, 2618, 2619: oled_data = 16'b1111111111111111;
    2620, 2621, 2622, 2623, 2624, 2625, 2626, 2627, 2628, 2629: oled_data = 16'b1111111111111111;
    2630, 2631, 2632, 2633, 2634, 2635, 2636, 2637, 2638, 2639: oled_data = 16'b1111111111111111;
    2640, 2641, 2642, 2643, 2644, 2645, 2646, 2647, 2648, 2649: oled_data = 16'b1111111111111111;
    2650, 2651, 2652, 2653, 2654, 2655, 2656, 2657, 2658, 2659: oled_data = 16'b1111111111111111;
    2685, 2686, 2687, 2688, 2689, 2690, 2691, 2692, 2693, 2694: oled_data = 16'b1111111111111111;
    2696, 2698, 2700, 2702, 2704, 2706, 2708, 2710, 2712, 2714: oled_data = 16'b1111111111111111;
    2716, 2718, 2720, 2722, 2724, 2728, 2730, 2732, 2734, 2736: oled_data = 16'b1111111111111111;
    2738, 2740, 2742, 2746, 2747, 2748, 2749, 2750, 2751, 2752: oled_data = 16'b1111111111111111;
    2753, 2754, 2781, 2782, 2783, 2784, 2785, 2786, 2787, 2845: oled_data = 16'b1111111111111111;
    2846, 2847, 2848, 2849, 2850, 2851, 2877, 2878, 2879, 2880: oled_data = 16'b1111111111111111;
    2881, 2943, 2944, 2945, 2946, 2947, 2973, 2974, 2975, 2976: oled_data = 16'b1111111111111111;
    2977, 3040, 3041, 3042, 3043, 3069, 3070, 3071, 3072, 3137: oled_data = 16'b1111111111111111;
    3138, 3139, 3165, 3166, 3167, 3233, 3234, 3235, 3261, 3262: oled_data = 16'b1111111111111111;
    3263, 3329, 3330, 3357, 3358, 3359, 3451, 3452, 3453, 3454: oled_data = 16'b1111111111111111;
    3455, 3520, 3546, 3579, 3583, 3598, 3641, 3642, 3675, 3679: oled_data = 16'b1111111111111111;
    3727, 3728, 3729, 3737, 3766, 3771, 3775, 3779, 3782, 3783: oled_data = 16'b1111111111111111;
    3784, 3790, 3820, 3867, 3871, 3880, 3886, 3955, 3958, 3977: oled_data = 16'b1111111111111111;
    4004, 4127, 4512, 4608, 4672, 4704, 4705, 4706, 4766, 4767: oled_data = 16'b1111111111111111;
    4768, 4769, 4770, 4771, 4772, 4800, 4801, 4802, 4803, 4860: oled_data = 16'b1111111111111111;
    4861, 4862, 4863, 4864, 4865, 4870, 4895, 4896, 4897, 4898: oled_data = 16'b1111111111111111;
    4899, 4900, 4901, 4902, 4903, 4904, 4905, 4907, 4908, 4909: oled_data = 16'b1111111111111111;
    4910, 4911, 4912, 4913, 4914, 4915, 4916, 4917, 4918, 4919: oled_data = 16'b1111111111111111;
    4920, 4921, 4922, 4923, 4924, 4925, 4926, 4927, 4928, 4929: oled_data = 16'b1111111111111111;
    4930, 4932, 4933, 4934, 4935, 4936, 4937, 4938, 4939, 4940: oled_data = 16'b1111111111111111;
    4942, 4943, 4944, 4945, 4946, 4947, 4949, 4950, 4951, 4952: oled_data = 16'b1111111111111111;
    4953, 4954, 4955, 4956, 4957, 4958, 4959, 4960, 4961, 4962: oled_data = 16'b1111111111111111;
    4963, 4964, 4965, 4966, 4990, 4991, 4992, 4993, 4994, 4995: oled_data = 16'b1111111111111111;
    4996, 4997, 4998, 4999, 5000, 5001, 5002, 5003, 5004, 5005: oled_data = 16'b1111111111111111;
    5006, 5007, 5008, 5009, 5010, 5011, 5012, 5013, 5014, 5015: oled_data = 16'b1111111111111111;
    5016, 5017, 5018, 5019, 5020, 5021, 5022, 5023, 5024, 5025: oled_data = 16'b1111111111111111;
    5026, 5027, 5028, 5029, 5030, 5031, 5032, 5033, 5034, 5035: oled_data = 16'b1111111111111111;
    5036, 5037, 5038, 5039, 5040, 5041, 5042, 5043, 5044, 5045: oled_data = 16'b1111111111111111;
    5046, 5047, 5048, 5049, 5050, 5051, 5052, 5053, 5054, 5055: oled_data = 16'b1111111111111111;
    5056, 5057, 5058, 5059, 5060, 5061, 5062, 5086, 5087, 5088: oled_data = 16'b1111111111111111;
    5089, 5090, 5091, 5092, 5093, 5094, 5095, 5096, 5097, 5098: oled_data = 16'b1111111111111111;
    5099, 5100, 5101, 5102, 5103, 5104, 5105, 5106, 5107, 5108: oled_data = 16'b1111111111111111;
    5109, 5110, 5111, 5112, 5113, 5114, 5115, 5116, 5117, 5118: oled_data = 16'b1111111111111111;
    5119, 5120, 5121, 5122, 5123, 5124, 5125, 5126, 5127, 5128: oled_data = 16'b1111111111111111;
    5129, 5130, 5131, 5132, 5133, 5134, 5135, 5136, 5137, 5138: oled_data = 16'b1111111111111111;
    5139, 5140, 5141, 5142, 5143, 5144, 5145, 5146, 5147, 5148: oled_data = 16'b1111111111111111;
    5149, 5150, 5151, 5152, 5153, 5154, 5155, 5156, 5157, 5158: oled_data = 16'b1111111111111111;
    5159, 5177, 5178, 5179, 5180, 5181, 5182, 5183, 5184, 5185: oled_data = 16'b1111111111111111;
    5186, 5187, 5188, 5189, 5190, 5191, 5192, 5193, 5194, 5195: oled_data = 16'b1111111111111111;
    5196, 5197, 5198, 5199, 5200, 5201, 5202, 5203, 5204, 5205: oled_data = 16'b1111111111111111;
    5206, 5207, 5208, 5209, 5210, 5211, 5212, 5213, 5214, 5215: oled_data = 16'b1111111111111111;
    5216, 5217, 5218, 5219, 5220, 5221, 5222, 5223, 5224, 5225: oled_data = 16'b1111111111111111;
    5226, 5227, 5228, 5229, 5230, 5231, 5232, 5233, 5234, 5235: oled_data = 16'b1111111111111111;
    5236, 5237, 5238, 5239, 5240, 5241, 5242, 5243, 5244, 5245: oled_data = 16'b1111111111111111;
    5246, 5247, 5248, 5249, 5250, 5251, 5252, 5253, 5254, 5255: oled_data = 16'b1111111111111111;
    5272, 5273, 5274, 5275, 5276, 5277, 5278, 5279, 5280, 5281: oled_data = 16'b1111111111111111;
    5282, 5283, 5284, 5285, 5286, 5287, 5288, 5289, 5290, 5291: oled_data = 16'b1111111111111111;
    5292, 5293, 5294, 5295, 5296, 5297, 5298, 5299, 5300, 5301: oled_data = 16'b1111111111111111;
    5302, 5303, 5304, 5305, 5306, 5307, 5308, 5309, 5310, 5311: oled_data = 16'b1111111111111111;
    5312, 5313, 5314, 5315, 5316, 5317, 5318, 5319, 5320, 5321: oled_data = 16'b1111111111111111;
    5322, 5323, 5324, 5325, 5326, 5327, 5328, 5329, 5330, 5331: oled_data = 16'b1111111111111111;
    5332, 5333, 5334, 5335, 5336, 5337, 5338, 5339, 5340, 5341: oled_data = 16'b1111111111111111;
    5342, 5343, 5344, 5345, 5346, 5347, 5348, 5349, 5350, 5351: oled_data = 16'b1111111111111111;
    5368, 5369, 5370, 5371, 5372, 5373, 5374, 5375, 5376, 5377: oled_data = 16'b1111111111111111;
    5378, 5379, 5380, 5381, 5382, 5383, 5384, 5385, 5386, 5387: oled_data = 16'b1111111111111111;
    5388, 5389, 5390, 5391, 5392, 5393, 5394, 5395, 5396, 5397: oled_data = 16'b1111111111111111;
    5398, 5399, 5400, 5401, 5402, 5403, 5404, 5405, 5406, 5407: oled_data = 16'b1111111111111111;
    5408, 5409, 5410, 5411, 5412, 5413, 5414, 5415, 5416, 5417: oled_data = 16'b1111111111111111;
    5418, 5419, 5420, 5421, 5422, 5423, 5424, 5425, 5426, 5427: oled_data = 16'b1111111111111111;
    5428, 5429, 5430, 5431, 5432, 5433, 5434, 5435, 5436, 5437: oled_data = 16'b1111111111111111;
    5438, 5439, 5440, 5441, 5442, 5443, 5444, 5445, 5446, 5447: oled_data = 16'b1111111111111111;
    5464, 5465, 5466, 5467, 5468, 5469, 5470, 5471, 5472, 5473: oled_data = 16'b1111111111111111;
    5474, 5475, 5476, 5477, 5478, 5479, 5480, 5481, 5482, 5483: oled_data = 16'b1111111111111111;
    5484, 5485, 5486, 5487, 5488, 5489, 5490, 5491, 5492, 5493: oled_data = 16'b1111111111111111;
    5494, 5495, 5496, 5497, 5498, 5499, 5500, 5501, 5502, 5503: oled_data = 16'b1111111111111111;
    5504, 5505, 5506, 5507, 5508, 5509, 5510, 5511, 5512, 5513: oled_data = 16'b1111111111111111;
    5514, 5515, 5516, 5517, 5518, 5519, 5520, 5521, 5522, 5523: oled_data = 16'b1111111111111111;
    5524, 5525, 5526, 5527, 5528, 5529, 5530, 5531, 5532, 5533: oled_data = 16'b1111111111111111;
    5534, 5535, 5536, 5537, 5538, 5539, 5540, 5542, 5560, 5561: oled_data = 16'b1111111111111111;
    5564, 5565, 5566, 5567, 5568, 5569, 5570, 5571, 5572, 5573: oled_data = 16'b1111111111111111;
    5574, 5575, 5576, 5577, 5578, 5579, 5580, 5581, 5582, 5583: oled_data = 16'b1111111111111111;
    5584, 5585, 5586, 5587, 5588, 5589, 5590, 5591, 5592, 5593: oled_data = 16'b1111111111111111;
    5594, 5595, 5596, 5597, 5598, 5599, 5600, 5601, 5602, 5603: oled_data = 16'b1111111111111111;
    5604, 5605, 5606, 5607, 5608, 5609, 5610, 5611, 5612, 5613: oled_data = 16'b1111111111111111;
    5614, 5615, 5616, 5617, 5618, 5619, 5620, 5621, 5622, 5623: oled_data = 16'b1111111111111111;
    5624, 5625, 5626, 5627, 5628, 5629, 5630, 5631, 5632, 5633: oled_data = 16'b1111111111111111;
    5634, 5635, 5664, 5665, 5666, 5667, 5668, 5669, 5670, 5671: oled_data = 16'b1111111111111111;
    5672, 5673, 5674, 5675, 5676, 5677, 5678, 5679, 5680, 5681: oled_data = 16'b1111111111111111;
    5682, 5683, 5684, 5685, 5686, 5687, 5688, 5689, 5690, 5691: oled_data = 16'b1111111111111111;
    5692, 5693, 5694, 5695, 5696, 5697, 5698, 5699, 5700, 5701: oled_data = 16'b1111111111111111;
    5702, 5703, 5704, 5705, 5706, 5707, 5708, 5709, 5710, 5711: oled_data = 16'b1111111111111111;
    5712, 5713, 5714, 5715, 5716, 5717, 5718, 5719, 5720, 5721: oled_data = 16'b1111111111111111;
    5722, 5723, 5724, 5725, 5726, 5727, 5728, 5729, 5730, 5760: oled_data = 16'b1111111111111111;
    5761, 5762, 5763, 5764, 5765, 5766, 5767, 5768, 5769, 5770: oled_data = 16'b1111111111111111;
    5771, 5772, 5773, 5774, 5775, 5776, 5777, 5778, 5779, 5780: oled_data = 16'b1111111111111111;
    5781, 5782, 5783, 5784, 5785, 5786, 5787, 5788, 5789, 5790: oled_data = 16'b1111111111111111;
    5791, 5792, 5793, 5794, 5795, 5796, 5797, 5798, 5799, 5800: oled_data = 16'b1111111111111111;
    5801, 5802, 5803, 5804, 5805, 5806, 5807, 5808, 5809, 5810: oled_data = 16'b1111111111111111;
    5811, 5812, 5813, 5814, 5815, 5816, 5817, 5818, 5819, 5820: oled_data = 16'b1111111111111111;
    5821, 5822, 5823, 5824, 5825, 5826, 5856, 5857, 5858, 5859: oled_data = 16'b1111111111111111;
    5860, 5861, 5862, 5863, 5864, 5865, 5866, 5867, 5868, 5869: oled_data = 16'b1111111111111111;
    5870, 5871, 5872, 5873, 5874, 5875, 5876, 5877, 5878, 5879: oled_data = 16'b1111111111111111;
    5880, 5881, 5882, 5883, 5884, 5885, 5886, 5887, 5888, 5889: oled_data = 16'b1111111111111111;
    5890, 5891, 5892, 5893, 5894, 5895, 5896, 5897, 5898, 5899: oled_data = 16'b1111111111111111;
    5900, 5901, 5902, 5903, 5904, 5905, 5906, 5907, 5908, 5909: oled_data = 16'b1111111111111111;
    5910, 5911, 5912, 5913, 5914, 5915, 5916, 5917, 5918, 5919: oled_data = 16'b1111111111111111;
    5920, 5921, 5922, 5923, 5952, 5953, 5954, 5955, 5956, 5957: oled_data = 16'b1111111111111111;
    5958, 5959, 5960, 5961, 5962, 5963, 5964, 5965, 5966, 5967: oled_data = 16'b1111111111111111;
    5968, 5969, 5970, 5971, 5972, 5973, 5974, 5975, 5976, 5977: oled_data = 16'b1111111111111111;
    5978, 5979, 5980, 5981, 5982, 5983, 5984, 5985, 5986, 5987: oled_data = 16'b1111111111111111;
    5988, 5989, 5990, 5991, 5992, 5993, 5994, 5995, 5996, 5997: oled_data = 16'b1111111111111111;
    5998, 5999, 6000, 6001, 6002, 6003, 6004, 6005, 6006, 6007: oled_data = 16'b1111111111111111;
    6008, 6009, 6010, 6011, 6012, 6013, 6014, 6015, 6016, 6017: oled_data = 16'b1111111111111111;
    6018, 6019, 6020, 6021, 6022, 6023, 6024, 6025, 6026, 6027: oled_data = 16'b1111111111111111;
    6028, 6029, 6030, 6031, 6032, 6033, 6034, 6035, 6036, 6037: oled_data = 16'b1111111111111111;
    6038, 6039, 6040, 6041, 6042, 6043, 6044, 6045, 6046, 6047: oled_data = 16'b1111111111111111;
    6048, 6049, 6050, 6051, 6052, 6053, 6054, 6055, 6056, 6057: oled_data = 16'b1111111111111111;
    6058, 6059, 6060, 6061, 6062, 6063, 6064, 6065, 6066, 6067: oled_data = 16'b1111111111111111;
    6068, 6069, 6070, 6071, 6072, 6073, 6074, 6075, 6076, 6077: oled_data = 16'b1111111111111111;
    6078, 6079, 6080, 6081, 6082, 6083, 6084, 6085, 6086, 6087: oled_data = 16'b1111111111111111;
    6088, 6089, 6090, 6091, 6092, 6093, 6094, 6095, 6096, 6097: oled_data = 16'b1111111111111111;
    6098, 6099, 6100, 6101, 6102, 6103, 6104, 6105, 6106, 6107: oled_data = 16'b1111111111111111;
    6108, 6109, 6110, 6111, 6112, 6113, 6114, 6115, 6116, 6117: oled_data = 16'b1111111111111111;
    6118, 6119, 6120, 6121, 6122, 6123, 6124, 6125, 6126, 6127: oled_data = 16'b1111111111111111;
    6128, 6129, 6130, 6131, 6132, 6133, 6134, 6135, 6136, 6137: oled_data = 16'b1111111111111111;
    6138, 6139, 6140, 6141, 6142, 6143: oled_data = 16'b1111111111111111;
    202, 241, 276, 782, 797, 1295, 1298, 2789, 2791, 2842: oled_data = 16'b1111011110111111;
    2883, 2941, 3073, 3135, 3264, 3328, 3500, 3685, 3957, 4128: oled_data = 16'b1111011110111111;
    4224, 4416, 4417, 4610, 4670, 4707, 4765, 4805, 4807, 4808: oled_data = 16'b1111011110111111;
    4810, 4812, 4814, 4815, 4817, 4818, 4820, 4821, 4825, 4827: oled_data = 16'b1111011110111111;
    4828, 4831, 4833, 4835, 4838, 4842, 4844, 4847, 4850, 4854: oled_data = 16'b1111011110111111;
    4856, 4858: oled_data = 16'b1111011110111111;
    211, 235, 258, 437, 521, 526, 537, 556, 656, 940: oled_data = 16'b1111111110111111;
    953, 1013, 1040, 1097, 1193, 1232, 1264, 1268, 1272, 1276: oled_data = 16'b1111111110111111;
    1280, 1294, 1307, 1311, 1315, 1319, 1333, 1719, 1816, 2695: oled_data = 16'b1111111110111111;
    2697, 2699, 2701, 2703, 2705, 2707, 2709, 2711, 2713, 2715: oled_data = 16'b1111111110111111;
    2717, 2719, 2721, 2723, 2725, 2727, 2729, 2731, 2733, 2735: oled_data = 16'b1111111110111111;
    2737, 2739, 2741, 2743, 2745, 2788, 2841, 2844, 2882, 2942: oled_data = 16'b1111111110111111;
    3039, 3168, 3232, 3356, 3360, 3425, 3589, 3690, 3694, 3776: oled_data = 16'b1111111110111111;
    3863, 3877, 3956, 3967, 4320, 4574, 4609, 4671, 4804, 4806: oled_data = 16'b1111111110111111;
    4809, 4811, 4822, 4824, 4829, 4832, 4836, 4839, 4841, 4845: oled_data = 16'b1111111110111111;
    4848, 4851, 4853, 4855, 4857, 4859, 4867, 4906, 4931, 4941: oled_data = 16'b1111111110111111;
    4948: oled_data = 16'b1111111110111111;
    212, 218, 226, 259, 265, 415, 435, 446, 495, 502: oled_data = 16'b1111011111111111;
    538, 549, 554, 561, 591, 687, 830, 857, 870, 922: oled_data = 16'b1111011111111111;
    938, 975, 1049, 1083, 1096, 1118, 1130, 1241, 1261, 1266: oled_data = 16'b1111011111111111;
    1286, 1292, 1304, 1327, 1331, 1335, 2726, 2744, 3823, 3912: oled_data = 16'b1111011111111111;
    3916, 4007, 5563: oled_data = 16'b1111011111111111;
    392, 2984, 2987, 2989, 2991, 2993, 2995, 2997, 3003, 3005: oled_data = 16'b1110010111111101;
    3007, 3009, 3011, 3013, 3015, 3017, 3019, 3021, 3023, 3025: oled_data = 16'b1110010111111101;
    3027, 3031, 3458, 3573, 3574, 3586, 3878, 4618, 4620, 4622: oled_data = 16'b1110010111111101;
    4624, 4631, 4641, 4644, 4646, 4654, 4656, 4658: oled_data = 16'b1110010111111101;
    393, 409, 456, 467: oled_data = 16'b1010010010111000;
    394: oled_data = 16'b1001110100111000;
    395, 403, 421, 432, 433, 450, 468, 1067: oled_data = 16'b1001110011111000;
    396, 404, 451: oled_data = 16'b1001010100111000;
    397: oled_data = 16'b1100111110111111;
    401, 1101: oled_data = 16'b1111111100111111;
    402: oled_data = 16'b1100010010111010;
    405, 452: oled_data = 16'b1100011101111110;
    408, 455, 466: oled_data = 16'b1111011000111110;
    410: oled_data = 16'b1011011010111100;
    412, 443: oled_data = 16'b1111111011111111;
    413: oled_data = 16'b1011110010111010;
    414, 469: oled_data = 16'b1001110111111010;
    416: oled_data = 16'b1111111010111110;
    417: oled_data = 16'b1010010001011000;
    418: oled_data = 16'b1010111011111100;
    420: oled_data = 16'b1110010110111101;
    422: oled_data = 16'b1011111101111110;
    426: oled_data = 16'b1101010100111011;
    427: oled_data = 16'b1001010101111001;
    428, 720: oled_data = 16'b1101011111111111;
    431: oled_data = 16'b1110110110111101;
    434: oled_data = 16'b1010011000111010;
    438: oled_data = 16'b1100110010111010;
    439: oled_data = 16'b1001010111111010;
    440, 511, 531, 616, 695, 742, 791, 838, 887, 934: oled_data = 16'b1101111111111111;
    983, 1030, 1079, 1126, 1175: oled_data = 16'b1101111111111111;
    444: oled_data = 16'b1011010010111001;
    445: oled_data = 16'b1001111001111011;
    448, 533, 617, 629, 725, 752, 821, 848, 917, 921: oled_data = 16'b1111111101111111;
    944, 1109, 1136, 1205: oled_data = 16'b1111111101111111;
    449: oled_data = 16'b1100010011111010;
    457: oled_data = 16'b1011011011111100;
    461: oled_data = 16'b1110010101111101;
    462: oled_data = 16'b1001010011111000;
    463: oled_data = 16'b1100111101111110;
    470, 542, 607, 638, 734, 820, 926, 1022, 1203, 1214: oled_data = 16'b1110111111111111;
    488: oled_data = 16'b1011101011011001;
    489: oled_data = 16'b0010100000001101;
    490, 854, 950: oled_data = 16'b0010100011001110;
    491, 635, 649, 1163: oled_data = 16'b0011100011001110;
    492: oled_data = 16'b0001100100001111;
    493: oled_data = 16'b0111011100111101;
    497, 923: oled_data = 16'b1111010110111110;
    498: oled_data = 16'b0110100001010011;
    499, 850: oled_data = 16'b0010100011001101;
    500, 547, 750: oled_data = 16'b0010000011001110;
    501, 548: oled_data = 16'b0110011001111011;
    504: oled_data = 16'b1110101111011110;
    505, 513, 552, 689, 736, 1073, 1081: oled_data = 16'b0011000000001101;
    506, 553: oled_data = 16'b0100110011110111;
    508: oled_data = 16'b1111110111111111;
    509: oled_data = 16'b0110100000010001;
    510: oled_data = 16'b0001001010010001;
    512, 608, 1088: oled_data = 16'b1111010010111110;
    514: oled_data = 16'b0010110011110111;
    516, 807: oled_data = 16'b1100001011011001;
    517: oled_data = 16'b0001100000001101;
    518: oled_data = 16'b0101111001111011;
    520, 1282: oled_data = 16'b1111011111111110;
    522: oled_data = 16'b1001000011010101;
    523: oled_data = 16'b0000100110001110;
    524: oled_data = 16'b1001011110111111;
    527: oled_data = 16'b1011101001011010;
    528, 977: oled_data = 16'b0011000001001110;
    529: oled_data = 16'b0011000001001101;
    530: oled_data = 16'b0010101101010100;
    534, 718, 910: oled_data = 16'b0111100001010011;
    535: oled_data = 16'b0001001000010000;
    536: oled_data = 16'b1010111110111111;
    539: oled_data = 16'b1110110101111110;
    540: oled_data = 16'b0100100000001110;
    541: oled_data = 16'b0001110000010101;
    544: oled_data = 16'b1111011001111110;
    545: oled_data = 16'b0110100011010011;
    546: oled_data = 16'b0010100010001101;
    551, 600, 743, 792, 839: oled_data = 16'b1111001111011110;
    555, 1256, 1259, 1274, 1297, 1313, 1330, 1805, 2588, 2684: oled_data = 16'b1111011110111110;
    2790, 2843, 2876, 2972, 2978, 3038, 3068, 3164, 3260, 3424: oled_data = 16'b1111011110111110;
    3481, 3547, 3594, 3630, 3725, 3767, 3781, 3963, 4101, 4102: oled_data = 16'b1111011110111110;
    4402, 4594, 4708, 4823, 4830, 4837, 4840, 4846, 4849, 4852: oled_data = 16'b1111011110111110;
    4869, 5085: oled_data = 16'b1111011110111110;
    557: oled_data = 16'b1011100111011001;
    558: oled_data = 16'b0001000001001101;
    559: oled_data = 16'b1000011010111100;
    562, 784: oled_data = 16'b1101001100011100;
    563: oled_data = 16'b0011100001001111;
    564, 777, 1201: oled_data = 16'b0011000010001101;
    565: oled_data = 16'b0010101010010010;
    566, 724, 1108: oled_data = 16'b1100011110111110;
    584, 612, 776, 872, 1064: oled_data = 16'b1100001100011010;
    585, 681, 709, 901, 969: oled_data = 16'b0010100010001110;
    586: oled_data = 16'b0110010111111010;
    587: oled_data = 16'b1110011101111110;
    588, 3576, 3613, 3651, 3939: oled_data = 16'b1101010010111100;
    589: oled_data = 16'b0101000011010000;
    590: oled_data = 16'b0100010011110111;
    592: oled_data = 16'b1110001101011100;
    593: oled_data = 16'b0100000100010000;
    594, 641: oled_data = 16'b0101010101111001;
    595, 642: oled_data = 16'b1101111101111110;
    596: oled_data = 16'b1101110010111101;
    597, 644: oled_data = 16'b0110000011010001;
    598, 645: oled_data = 16'b0011110000010110;
    599, 646, 1087, 1183, 1222: oled_data = 16'b1110011111111111;
    601, 697, 744, 832, 840, 936, 985, 1032: oled_data = 16'b0011100000001110;
    602, 698, 841: oled_data = 16'b0101110101111000;
    603: oled_data = 16'b1110111010111111;
    604: oled_data = 16'b1010001111011001;
    605: oled_data = 16'b0110101001010101;
    606: oled_data = 16'b0110110010110111;
    609, 685, 793, 801, 889, 993: oled_data = 16'b0100000000001110;
    610, 994: oled_data = 16'b0011110100110111;
    613, 1200: oled_data = 16'b0011100010001110;
    614, 906: oled_data = 16'b0011100011001101;
    615, 1213: oled_data = 16'b0011010001010110;
    618: oled_data = 16'b1001100101010110;
    619, 811: oled_data = 16'b0001100111001111;
    620, 716, 812, 908, 1100: oled_data = 16'b1001111111111111;
    621, 909: oled_data = 16'b1111111010111111;
    622, 4049, 4152: oled_data = 16'b1000100100010101;
    623: oled_data = 16'b0011001011010010;
    624: oled_data = 16'b1011011011111101;
    625, 2889, 2891, 2893, 2894, 2897, 2899, 2900, 2902, 2903: oled_data = 16'b1110111010111110;
    2905, 2907, 2909, 2911, 2913, 2915, 2917, 2919, 2921, 2923: oled_data = 16'b1110111010111110;
    2925, 2927, 2929, 2931, 2933, 2935, 3075, 3133, 3881, 4515: oled_data = 16'b1110111010111110;
    4613, 4667: oled_data = 16'b1110111010111110;
    626: oled_data = 16'b1001100110010111;
    627, 808: oled_data = 16'b0001100100001110;
    628: oled_data = 16'b1001011100111101;
    630, 4379: oled_data = 16'b0111100100010100;
    631: oled_data = 16'b0011000011001101;
    632: oled_data = 16'b0010100101001110;
    633, 1190: oled_data = 16'b0111011010111100;
    634, 1160: oled_data = 16'b1100001101011010;
    636, 789, 836: oled_data = 16'b0011100010001101;
    637: oled_data = 16'b0011010000010110;
    639: oled_data = 16'b1110010001011100;
    640: oled_data = 16'b0100000011010000;
    643, 3267, 3325, 3421, 4285, 4420: oled_data = 16'b1101110101111101;
    647, 696, 888, 935, 1127: oled_data = 16'b1111001111011101;
    648, 905, 1224: oled_data = 16'b0100000001001111;
    650: oled_data = 16'b0010101100010010;
    651: oled_data = 16'b1101011000111111;
    652, 1206: oled_data = 16'b1000100100010100;
    653: oled_data = 16'b0011000100001101;
    654: oled_data = 16'b0010100100001111;
    655, 847: oled_data = 16'b1000011011111011;
    657: oled_data = 16'b1010000101010111;
    658: oled_data = 16'b0010101001010000;
    659: oled_data = 16'b1010011010111101;
    660, 2886, 2887, 2888, 2890, 2892, 2895, 2898, 2904, 2908: oled_data = 16'b1110111011111110;
    2910, 2914, 2916, 2918, 2920, 2922, 2926, 2928, 2930, 2932: oled_data = 16'b1110111011111110;
    2934, 2936, 2937, 2980, 3036, 3170, 3230, 3457, 3479, 3483: oled_data = 16'b1110111011111110;
    3502, 3553, 3578, 3649, 3689, 3745, 3841, 3937, 4033, 4418: oled_data = 16'b1110111011111110;
    4573, 4713, 4714, 4715, 4716, 4717, 4718, 4719, 4720, 4721: oled_data = 16'b1110111011111110;
    4722, 4723, 4724, 4725, 4726, 4727, 4728, 4729, 4730, 4731: oled_data = 16'b1110111011111110;
    4732, 4733, 4734, 4735, 4736, 4737, 4738, 4739, 4740, 4741: oled_data = 16'b1110111011111110;
    4742, 4743, 4744, 4745, 4746, 4747, 4748, 4749, 4750, 4751: oled_data = 16'b1110111011111110;
    4752, 4753, 4754, 4755, 4756, 4757, 4758, 4759, 4760: oled_data = 16'b1110111011111110;
    661, 3873: oled_data = 16'b1011001011011010;
    662: oled_data = 16'b0011000101010000;
    663, 1239: oled_data = 16'b1000011001111011;
    680, 900, 968: oled_data = 16'b1100001100011001;
    682, 1094: oled_data = 16'b0110011010111100;
    684: oled_data = 16'b1111010100111110;
    686: oled_data = 16'b0010110010110110;
    688, 976, 1072: oled_data = 16'b1101101011011011;
    690: oled_data = 16'b0100110111111010;
    692: oled_data = 16'b1111010100111111;
    693, 981, 1028, 1077: oled_data = 16'b0110000000010000;
    694: oled_data = 16'b0001101111010100;
    699: oled_data = 16'b1101001101011101;
    700: oled_data = 16'b0010000000001101;
    701: oled_data = 16'b0110111000111010;
    704, 896, 904: oled_data = 16'b1110110011111110;
    705, 897: oled_data = 16'b0100000000001101;
    706, 898: oled_data = 16'b0011010100111000;
    708, 996: oled_data = 16'b1100101011011001;
    710, 1069: oled_data = 16'b0101101101010101;
    711, 747: oled_data = 16'b0111001011010110;
    712: oled_data = 16'b0111010010110110;
    713, 816: oled_data = 16'b1100111101111111;
    714: oled_data = 16'b1010000101010110;
    715: oled_data = 16'b0001000111001111;
    717, 813, 1005: oled_data = 16'b1111111001111111;
    719: oled_data = 16'b0010001010010001;
    722: oled_data = 16'b1110010100111100;
    723: oled_data = 16'b1001010010110111;
    726: oled_data = 16'b1000000011010011;
    727: oled_data = 16'b0010100111001111;
    728: oled_data = 16'b0111001110010110;
    729: oled_data = 16'b0110101100010110;
    730: oled_data = 16'b0110101101010110;
    731, 748: oled_data = 16'b0111001100010110;
    732: oled_data = 16'b0101000001001110;
    733, 1117: oled_data = 16'b0010010000010110;
    735, 927, 1119: oled_data = 16'b1101101111011011;
    737, 978, 1025: oled_data = 16'b0101010111111010;
    739, 1123: oled_data = 16'b1111010111111111;
    740: oled_data = 16'b0101100000010000;
    741, 1078: oled_data = 16'b0010001110010100;
    745: oled_data = 16'b0100101100010010;
    746: oled_data = 16'b1000001011010111;
    749, 3995: oled_data = 16'b1000000110010011;
    751, 943, 1039, 1135: oled_data = 16'b1000011011111100;
    753, 1041, 1137: oled_data = 16'b1001000010010101;
    754, 1138: oled_data = 16'b0001100110001111;
    755: oled_data = 16'b1011011111111110;
    757: oled_data = 16'b1100101010011010;
    758, 1065: oled_data = 16'b0010100001001101;
    759: oled_data = 16'b0111011000111011;
    774, 1131, 1284, 2780, 3777, 4209, 4498, 4513, 4813, 4816: oled_data = 16'b1111111110111110;
    4819, 4826, 4834, 4843, 5541, 5562: oled_data = 16'b1111111110111110;
    778, 786, 787, 788, 834, 851, 852: oled_data = 16'b0011100101001111;
    779: oled_data = 16'b0100000101001111;
    780: oled_data = 16'b0010100110010000;
    781: oled_data = 16'b0111011010111101;
    785: oled_data = 16'b0100000001001110;
    790, 933: oled_data = 16'b0010101110010101;
    794: oled_data = 16'b0011100100001110;
    795: oled_data = 16'b0011001010010010;
    796: oled_data = 16'b1010111100111101;
    800, 992: oled_data = 16'b1110110010111110;
    802: oled_data = 16'b0011110011110111;
    804: oled_data = 16'b1100101100011010;
    805: oled_data = 16'b0010000010001101;
    806: oled_data = 16'b0111011011111101;
    809: oled_data = 16'b0111111001111101;
    810: oled_data = 16'b1001100101010101;
    814: oled_data = 16'b1000000001010011;
    815: oled_data = 16'b0010001011010001;
    817, 3596, 3687: oled_data = 16'b1101110111111100;
    818: oled_data = 16'b1011111000111100;
    819: oled_data = 16'b1100011010111100;
    822, 918, 1014, 1110: oled_data = 16'b1000000010010011;
    823: oled_data = 16'b0001101011010010;
    824: oled_data = 16'b1011011011111111;
    825: oled_data = 16'b1000100010010010;
    826: oled_data = 16'b0010010001010100;
    827: oled_data = 16'b1101010111111111;
    828, 1124: oled_data = 16'b0101100000001111;
    829: oled_data = 16'b0010010001010101;
    831: oled_data = 16'b1101101111011100;
    833: oled_data = 16'b0011100101001110;
    835: oled_data = 16'b0011100110001111;
    837, 886: oled_data = 16'b0010101111010101;
    842: oled_data = 16'b1110010000011101;
    843, 873: oled_data = 16'b0011000010001110;
    844: oled_data = 16'b1000011001111100;
    845: oled_data = 16'b1101001010011011;
    846, 942, 997, 1038: oled_data = 16'b0010000010001110;
    849, 945: oled_data = 16'b1001000011010110;
    853, 1189: oled_data = 16'b0011100100001111;
    855, 1047, 1143: oled_data = 16'b0111111001111011;
    874: oled_data = 16'b0100101101010100;
    875: oled_data = 16'b1001001111010101;
    876: oled_data = 16'b0111101011010101;
    877: oled_data = 16'b0110110000010111;
    878: oled_data = 16'b1010111010111011;
    880: oled_data = 16'b1101101100011100;
    881, 928: oled_data = 16'b0011100001001110;
    882, 929: oled_data = 16'b0100001100010011;
    883, 930: oled_data = 16'b1000110000010110;
    884: oled_data = 16'b1000101011010110;
    885, 932: oled_data = 16'b0100100001001110;
    890: oled_data = 16'b0100101011010010;
    891: oled_data = 16'b0111101011010111;
    892: oled_data = 16'b0111110001010111;
    893: oled_data = 16'b1100011100111100;
    902: oled_data = 16'b0110111001111011;
    907, 1003: oled_data = 16'b0010000111010000;
    911: oled_data = 16'b0010101100010001;
    912: oled_data = 16'b1100110101111111;
    913, 3413, 3415, 3416, 4135: oled_data = 16'b0110100001010010;
    914: oled_data = 16'b0010000011001101;
    915: oled_data = 16'b0010000100001111;
    916: oled_data = 16'b1000111100111100;
    919, 1015: oled_data = 16'b0001101010010001;
    920, 1043: oled_data = 16'b1011011110111111;
    924: oled_data = 16'b0101000000001111;
    925: oled_data = 16'b0010110000010110;
    931: oled_data = 16'b1000101100010110;
    937, 1129: oled_data = 16'b0101010100110111;
    939, 1257, 1260, 1277, 1290, 1296, 1302, 1308, 1316, 1320: oled_data = 16'b1111011101111110;
    1329, 1809, 2491, 2792, 2794, 2796, 2798, 2800, 2802, 2804: oled_data = 16'b1111011101111110;
    2806, 2808, 2810, 2812, 2814, 2816, 2818, 2820, 2822, 2824: oled_data = 16'b1111011101111110;
    2826, 2828, 2830, 2832, 2834, 2836, 2838, 2840, 2884, 3037: oled_data = 16'b1111011101111110;
    3169, 3327, 3476, 3478, 3484, 3485, 3488, 3489, 3494, 3495: oled_data = 16'b1111011101111110;
    3496, 3503, 3587, 3648, 3683, 3764, 3785, 3876, 3917, 3936: oled_data = 16'b1111011101111110;
    3973, 3982, 4611: oled_data = 16'b1111011101111110;
    941: oled_data = 16'b1100001000011001;
    946: oled_data = 16'b0010100101001101;
    947: oled_data = 16'b0111001111010110;
    948: oled_data = 16'b1001001111010110;
    949, 3611: oled_data = 16'b0111100110010100;
    951: oled_data = 16'b0111111000111011;
    970: oled_data = 16'b0110111011111100;
    972: oled_data = 16'b1111010101111110;
    973: oled_data = 16'b0011100000001100;
    974: oled_data = 16'b0001010000010101;
    980: oled_data = 16'b1111110100111111;
    982, 1029: oled_data = 16'b0010001111010100;
    984: oled_data = 16'b1111001110011110;
    986: oled_data = 16'b0101110110111000;
    987: oled_data = 16'b1101101111011101;
    988, 1024, 1120: oled_data = 16'b0011000000001110;
    989: oled_data = 16'b0110010100111001;
    990, 1321: oled_data = 16'b1110111110111111;
    998: oled_data = 16'b0110111010111100;
    1000: oled_data = 16'b1111011010111110;
    1001: oled_data = 16'b1011010010111010;
    1002: oled_data = 16'b0110100101010010;
    1004: oled_data = 16'b1001011111111110;
    1006: oled_data = 16'b0111100000010011;
    1007: oled_data = 16'b0001101010010000;
    1008: oled_data = 16'b1101011110111111;
    1009, 2985, 2992, 2998, 3000, 3008, 3020, 3032, 3614, 4626: oled_data = 16'b1110010111111110;
    4628, 4634, 4636, 4638, 4649, 4651, 4661: oled_data = 16'b1110010111111110;
    1010: oled_data = 16'b1001000110010101;
    1011: oled_data = 16'b0001100001001101;
    1012: oled_data = 16'b1000011100111101;
    1016, 1112, 1208: oled_data = 16'b1011011111111111;
    1019, 1115, 1211: oled_data = 16'b1111010110111111;
    1020, 1116: oled_data = 16'b0101000000001110;
    1021: oled_data = 16'b0010110001010110;
    1023: oled_data = 16'b1110001111011011;
    1027, 1180, 1219: oled_data = 16'b1111111000111111;
    1031, 1080: oled_data = 16'b1111101111011110;
    1033: oled_data = 16'b0101110100111000;
    1037: oled_data = 16'b1100001001011001;
    1042: oled_data = 16'b0010000111001111;
    1045: oled_data = 16'b1101001011011010;
    1046: oled_data = 16'b0010100001001110;
    1066: oled_data = 16'b0100101111010101;
    1068: oled_data = 16'b1000101101010111;
    1070: oled_data = 16'b1000111000111011;
    1074: oled_data = 16'b0100110110111001;
    1076, 1184: oled_data = 16'b1111010011111110;
    1082: oled_data = 16'b0101010011111000;
    1084: oled_data = 16'b1111110110111110;
    1085: oled_data = 16'b0111000010010010;
    1086: oled_data = 16'b0010101100010011;
    1089, 1128: oled_data = 16'b0011100000001101;
    1090: oled_data = 16'b0011010011110111;
    1092: oled_data = 16'b1100001011011010;
    1093, 1142: oled_data = 16'b0010000001001101;
    1098: oled_data = 16'b1001100100010101;
    1099: oled_data = 16'b0001000110001111;
    1102, 3654, 3750, 3898: oled_data = 16'b1011001110011001;
    1103: oled_data = 16'b0110101010010101;
    1104: oled_data = 16'b1000010010110111;
    1105: oled_data = 16'b1010110011111000;
    1106: oled_data = 16'b0111101010010111;
    1107: oled_data = 16'b0110101111010101;
    1111: oled_data = 16'b0001101001010001;
    1121: oled_data = 16'b0100110111111001;
    1125: oled_data = 16'b0010001110010101;
    1133: oled_data = 16'b1100001000011010;
    1134: oled_data = 16'b0001100010001101;
    1139, 1235: oled_data = 16'b1011011110111110;
    1141, 1229: oled_data = 16'b1100001010011010;
    1161, 1169: oled_data = 16'b0100000011001111;
    1162: oled_data = 16'b0100100100001110;
    1164: oled_data = 16'b0010000101001111;
    1165: oled_data = 16'b1000111110111110;
    1168: oled_data = 16'b1101101101011100;
    1170, 1217: oled_data = 16'b0101110111111010;
    1172: oled_data = 16'b1111110101111111;
    1173: oled_data = 16'b0110100001010001;
    1174, 1221: oled_data = 16'b0011010000010101;
    1176, 1223: oled_data = 16'b1111010000011110;
    1177: oled_data = 16'b0100100001001111;
    1178: oled_data = 16'b0110010101111000;
    1181, 4137, 4139: oled_data = 16'b0111100010010011;
    1182: oled_data = 16'b0011001101010011;
    1185: oled_data = 16'b0100100010001111;
    1186: oled_data = 16'b0100010100111000;
    1188: oled_data = 16'b1100101101011010;
    1192, 1808, 1902, 1914, 2468, 2755, 3136, 3243, 3250, 3632: oled_data = 16'b1111111111111110;
    4491, 4690, 4786, 4866, 4868: oled_data = 16'b1111111111111110;
    1194: oled_data = 16'b1010000110010110;
    1195: oled_data = 16'b0010001001010000;
    1196: oled_data = 16'b1010011111111111;
    1199: oled_data = 16'b1101001100011011;
    1202: oled_data = 16'b0011001111010100;
    1207: oled_data = 16'b0010101011010010;
    1212: oled_data = 16'b0110000010010000;
    1215: oled_data = 16'b1110010000011100;
    1216: oled_data = 16'b0011100010001111;
    1220: oled_data = 16'b0110100010010001;
    1225: oled_data = 16'b0110010100111000;
    1230: oled_data = 16'b0011000100001111;
    1231: oled_data = 16'b1000111011111100;
    1233: oled_data = 16'b1001100100010110;
    1234: oled_data = 16'b0010101000010000;
    1237: oled_data = 16'b1101001011011011;
    1238: oled_data = 16'b0011000011001111;
    1258, 1270, 1278, 1291, 1303, 1309, 1317: oled_data = 16'b1110111110111110;
    1265, 1269, 1273, 1281, 1285, 1312, 1326, 1334: oled_data = 16'b1110111101111110;
    1325, 4764: oled_data = 16'b1111111101111110;
    1705, 5463: oled_data = 16'b1110011100111011;
    1706, 1715, 1716, 1717, 3548, 3631, 3822, 3824, 5367, 5747: oled_data = 16'b1110011011111011;
    1707, 5827: oled_data = 16'b1101111010111010;
    1708, 1714, 1999, 3331, 3551, 3629, 3634, 3730, 3921, 4100: oled_data = 16'b1110111101111101;
    4113, 4306, 5951: oled_data = 16'b1110111101111101;
    1718, 3550, 3918, 5737: oled_data = 16'b1101111011111010;
    1800, 5081, 5543: oled_data = 16'b1101111010111001;
    1801: oled_data = 16'b1001101110001011;
    1802, 1812, 4606: oled_data = 16'b1001001101001001;
    1803, 1911, 2761, 4315: oled_data = 16'b0111001010000110;
    1804, 2181, 2298: oled_data = 16'b1010010001010000;
    1810: oled_data = 16'b1011110100110001;
    1811, 1991, 4872, 4968: oled_data = 16'b1000101100001000;
    1813: oled_data = 16'b1001001100001001;
    1814, 3544: oled_data = 16'b0111001010000111;
    1815, 3999: oled_data = 16'b1100111001110111;
    1895, 3355, 3640, 3738, 4871, 5083, 5640: oled_data = 16'b1101011001111000;
    1896, 4986: oled_data = 16'b1001001101001010;
    1897, 2199, 2295, 2391, 4123: oled_data = 16'b1110110100101010;
    1898, 2383: oled_data = 16'b1110110100101001;
    1899, 2284: oled_data = 16'b1101110001000110;
    1900: oled_data = 16'b1001001100000100;
    1901: oled_data = 16'b1000101110001110;
    1905, 5734: oled_data = 16'b1000001110001101;
    1906: oled_data = 16'b1010101110001000;
    1907, 2375: oled_data = 16'b1111110110101011;
    1908: oled_data = 16'b1110110101101001;
    1909: oled_data = 16'b1110010011101000;
    1910, 3637, 5358, 5454, 5461, 5550, 5557, 5646: oled_data = 16'b1100110000000101;
    1912, 4894, 5660: oled_data = 16'b1100010111110111;
    1990, 3450: oled_data = 16'b1011110110110110;
    1992, 4796: oled_data = 16'b1110010100101010;
    1993, 4971: oled_data = 16'b1111011011110111;
    1994: oled_data = 16'b1110111000110011;
    1995: oled_data = 16'b1110110100101011;
    1996, 4886, 4887: oled_data = 16'b1101010001000101;
    1997, 2182, 2374, 2867: oled_data = 16'b1010101110000110;
    1998, 2394, 3839: oled_data = 16'b1010010001001111;
    2000, 4676: oled_data = 16'b1010010000001111;
    2001: oled_data = 16'b1100010000001000;
    2002, 2574, 3539: oled_data = 16'b1111011000110001;
    2003: oled_data = 16'b1111111101111010;
    2004: oled_data = 16'b1111011010110111;
    2005, 2102, 3348: oled_data = 16'b1110010110110000;
    2006, 5173: oled_data = 16'b1110010011100111;
    2007, 4212, 5259: oled_data = 16'b1100101111000101;
    2008: oled_data = 16'b1000001011000111;
    2009, 4799, 5841: oled_data = 16'b1011010101110100;
    2085, 3736: oled_data = 16'b1100010111110110;
    2086, 5065: oled_data = 16'b1010101111001010;
    2087: oled_data = 16'b1100110010101010;
    2088: oled_data = 16'b1111111011110110;
    2089, 3242, 3338, 3346, 3919, 4204, 4206, 4302, 4395, 4587: oled_data = 16'b1111111110111101;
    4683, 4882, 4972, 4976: oled_data = 16'b1111111110111101;
    2090: oled_data = 16'b1110111001110110;
    2091, 2764, 4596: oled_data = 16'b1110110101101100;
    2092, 5076, 5165, 5166: oled_data = 16'b1110010010100110;
    2093, 2285, 2778, 2874: oled_data = 16'b1011101110000101;
    2094, 3259, 4775, 5353: oled_data = 16'b1000101101001011;
    2095, 4108, 4304, 4495, 4592, 4974, 5736: oled_data = 16'b1111011101111101;
    2096, 3625, 4410, 5751: oled_data = 16'b0110101010001000;
    2097, 5162: oled_data = 16'b1100110001000111;
    2098, 2477, 2953: oled_data = 16'b1111111011110100;
    2100, 3147, 3151, 3248, 3343, 3345, 3434, 4016, 4110, 4111: oled_data = 16'b1111111110111100;
    4205, 4208, 4303, 4305, 4399, 4400, 4493, 4494, 4496, 4497: oled_data = 16'b1111111110111100;
    4588, 4590, 4591, 4593, 4684, 4687, 4688, 4781, 4878, 4879: oled_data = 16'b1111111110111100;
    4973: oled_data = 16'b1111111110111100;
    2101, 2185, 2293, 5458: oled_data = 16'b1111011011111001;
    2103: oled_data = 16'b1110010100101000;
    2104: oled_data = 16'b1011101110000100;
    2105, 4702: oled_data = 16'b1001001101001000;
    2106: oled_data = 16'b1010110100110100;
    2183, 2773, 5071: oled_data = 16'b1111111001101111;
    2184, 3344, 3821, 3825, 4223, 4397, 4975, 5063: oled_data = 16'b1111011110111101;
    2186: oled_data = 16'b1110010111110101;
    2187, 3161: oled_data = 16'b1110010101101100;
    2188, 2392, 5164, 5261: oled_data = 16'b1110010010100101;
    2189, 4579: oled_data = 16'b1011101111000110;
    2190, 4510, 5161, 5449: oled_data = 16'b1000001100001010;
    2191: oled_data = 16'b1011010100110011;
    2192: oled_data = 16'b0110101010001001;
    2193, 4309: oled_data = 16'b1101010001000111;
    2194, 4595: oled_data = 16'b1111111001110010;
    2195, 3049, 3144, 3535, 3537, 5452: oled_data = 16'b1110111011111001;
    2196, 4008: oled_data = 16'b1111011011111010;
    2197, 3050, 3153, 4685, 4782, 4784, 4876: oled_data = 16'b1111011110111100;
    2198: oled_data = 16'b1110110111110101;
    2200, 5163: oled_data = 16'b1110110011100110;
    2201: oled_data = 16'b1001101011000100;
    2202, 4798: oled_data = 16'b1000101110001101;
    2277: oled_data = 16'b1010110010110001;
    2278, 4287: oled_data = 16'b1010101110000111;
    2279, 2862, 3446: oled_data = 16'b1111111000101110;
    2280: oled_data = 16'b1111011010111001;
    2281: oled_data = 16'b1110110111110000;
    2282, 4388: oled_data = 16'b1110110110110000;
    2283, 2388, 2955, 4413: oled_data = 16'b1111010101101011;
    2286: oled_data = 16'b1010101110001001;
    2287: oled_data = 16'b1010001110000111;
    2288, 4121: oled_data = 16'b1001001011000111;
    2289: oled_data = 16'b1101110010101001;
    2290: oled_data = 16'b1111010110101101;
    2291: oled_data = 16'b1110110110101111;
    2292, 4200, 4389: oled_data = 16'b1110110111110010;
    2294, 3913: oled_data = 16'b1110010111110100;
    2296: oled_data = 16'b1101110010100101;
    2297, 2393, 2489: oled_data = 16'b1010001101000101;
    2373, 3426: oled_data = 16'b1010010001010001;
    2376, 2390, 4197: oled_data = 16'b1110110110110001;
    2377, 3541, 4696, 4885, 4970, 4978, 4979: oled_data = 16'b1111010101101010;
    2378, 2387: oled_data = 16'b1111010101101000;
    2379, 4019, 4884, 5645: oled_data = 16'b1111010100100111;
    2380: oled_data = 16'b1101010000001000;
    2381, 4581, 5364: oled_data = 16'b1100110000001001;
    2382, 2859: oled_data = 16'b1111110111101011;
    2384, 3062: oled_data = 16'b1100001101000110;
    2385, 3836, 4873, 5066, 5170: oled_data = 16'b1110110011101000;
    2386, 2471, 2474, 2481, 2482, 2566, 2579, 2580, 2582, 2665: oled_data = 16'b1111110110101010;
    2674, 2863, 2871, 3445, 3742, 5073: oled_data = 16'b1111110110101010;
    2389, 4888, 5460: oled_data = 16'b1110010111110010;
    2469, 5839: oled_data = 16'b1001001111001110;
    2470, 4577: oled_data = 16'b1001101101000110;
    2472: oled_data = 16'b1111010110101010;
    2473, 2483, 2485, 2568, 2578, 2581, 2583, 2677, 2678, 3827: oled_data = 16'b1111110101101001;
    3830, 4312, 5549: oled_data = 16'b1111110101101001;
    2475, 2585, 4700: oled_data = 16'b1100101110000110;
    2476, 2572, 2668: oled_data = 16'b1101010001001011;
    2478: oled_data = 16'b1111010111110001;
    2479, 3157, 4412, 4777, 5556: oled_data = 16'b1011101101000110;
    2480, 2956, 2957, 2958, 4316: oled_data = 16'b1111010100101010;
    2484, 2567, 2774: oled_data = 16'b1111110101101010;
    2486, 2487, 2584, 2675, 2679, 2775, 2872: oled_data = 16'b1111010101101001;
    2488, 2873, 3732, 4980: oled_data = 16'b1110110011100111;
    2490: oled_data = 16'b1001110000001111;
    2564: oled_data = 16'b1001110000001110;
    2565, 3528, 4313: oled_data = 16'b1100010001001001;
    2569, 2676, 4598, 4599: oled_data = 16'b1111010100101000;
    2570, 4977: oled_data = 16'b1111111001110001;
    2571: oled_data = 16'b1100010000001010;
    2573: oled_data = 16'b1111111100110101;
    2575, 2671, 3063, 5547: oled_data = 16'b1011101100000110;
    2576, 2672: oled_data = 16'b1111011000110010;
    2577, 2860, 5067: oled_data = 16'b1111110111101100;
    2586: oled_data = 16'b1000001000000100;
    2587: oled_data = 16'b0111101101001011;
    2660, 2852: oled_data = 16'b1001001110001101;
    2661, 3045, 3543: oled_data = 16'b1010001011000110;
    2662, 2966, 3350: oled_data = 16'b1101110001000111;
    2663: oled_data = 16'b1111110101101000;
    2664: oled_data = 16'b1111110111101010;
    2666, 4499: oled_data = 16'b1111111010110010;
    2667: oled_data = 16'b1100001111001001;
    2669, 2765, 3432, 3838: oled_data = 16'b1111111011110101;
    2670, 3922: oled_data = 16'b1110111000110001;
    2673: oled_data = 16'b1111111000101101;
    2680, 4291: oled_data = 16'b1100101111000110;
    2681, 4117: oled_data = 16'b1100001110000101;
    2682: oled_data = 16'b1010101101000100;
    2683: oled_data = 16'b1000101101001100;
    2756, 2948, 3044: oled_data = 16'b1001001111001101;
    2757: oled_data = 16'b1011001101000110;
    2758: oled_data = 16'b1111010101101100;
    2759: oled_data = 16'b1101010101101101;
    2760: oled_data = 16'b0110101010000110;
    2762: oled_data = 16'b1101110111110001;
    2763: oled_data = 16'b1110110100101100;
    2766, 4114, 4691, 4883: oled_data = 16'b1111011001110010;
    2767, 2868, 5554: oled_data = 16'b1110010010101001;
    2768: oled_data = 16'b1111111010110011;
    2769: oled_data = 16'b1001101111001010;
    2770: oled_data = 16'b0101101001000101;
    2771: oled_data = 16'b1011010000000111;
    2772: oled_data = 16'b1111111000101100;
    2776, 4120: oled_data = 16'b1110010001000111;
    2777, 3733: oled_data = 16'b1101010001000110;
    2779: oled_data = 16'b1001001111001100;
    2793, 2795, 2797, 2799, 2801, 2803, 2805, 2807, 2809, 2811: oled_data = 16'b1111011101111111;
    2813, 2815, 2817, 2819, 2821, 2823, 2825, 2827, 2829, 2831: oled_data = 16'b1111011101111111;
    2833, 2835, 2837, 2839, 2940, 3134, 3231, 3456, 3477, 3490: oled_data = 16'b1111011101111111;
    3552, 3571, 3744, 3778, 3840, 4032, 4514, 4669, 4709, 4763: oled_data = 16'b1111011101111111;
    2853: oled_data = 16'b1100110010101000;
    2854, 2864, 2960: oled_data = 16'b1111110111101101;
    2855: oled_data = 16'b1011110001001011;
    2856: oled_data = 16'b0111101011000110;
    2857: oled_data = 16'b0111101101001010;
    2858: oled_data = 16'b1110010110101110;
    2861, 5069, 5070: oled_data = 16'b1111111000101111;
    2865: oled_data = 16'b1001110000001100;
    2866: oled_data = 16'b0110101011000111;
    2869: oled_data = 16'b1101110011101101;
    2870, 3837, 4795, 5074: oled_data = 16'b1111110110101001;
    2875, 3140, 4774: oled_data = 16'b1001001110001100;
    2885, 2939, 3074, 3265, 3423, 3482, 3497, 3501, 3504, 3519: oled_data = 16'b1111011100111110;
    3666, 3667, 3684, 3763, 3765, 3780, 3978, 4225, 4321, 4710: oled_data = 16'b1111011100111110;
    4761, 4762: oled_data = 16'b1111011100111110;
    2896, 4322: oled_data = 16'b1110011010111110;
    2901, 2906, 2912, 2924: oled_data = 16'b1110011011111110;
    2938, 3686, 3972, 4129, 4712: oled_data = 16'b1111011011111110;
    2949, 4580: oled_data = 16'b1011101111001000;
    2950: oled_data = 16'b1101001111000111;
    2951: oled_data = 16'b1100101110000111;
    2952: oled_data = 16'b1111110110101100;
    2954: oled_data = 16'b1111111000110000;
    2959, 4695: oled_data = 16'b1111010111101110;
    2961: oled_data = 16'b1111111010110100;
    2962: oled_data = 16'b1111111001110000;
    2963: oled_data = 16'b1101110000000111;
    2964: oled_data = 16'b1011001011000110;
    2965, 3064: oled_data = 16'b1011101101000111;
    2967, 4681: oled_data = 16'b1110010010101000;
    2968, 5169: oled_data = 16'b1101110010100111;
    2969: oled_data = 16'b1101010000000110;
    2970: oled_data = 16'b1010001101000100;
    2971, 4029, 5655: oled_data = 16'b1000101110001100;
    2979, 4478: oled_data = 16'b1111011100111111;
    2981, 3035, 3266, 3326, 3875, 4666: oled_data = 16'b1110011001111110;
    2982, 2983, 3034, 3422, 3580, 4615, 4617, 4619, 4621, 4623: oled_data = 16'b1110011000111110;
    4625, 4630, 4632, 4640, 4642, 4643, 4645, 4647, 4653, 4655: oled_data = 16'b1110011000111110;
    4657, 4659, 4664: oled_data = 16'b1110011000111110;
    2986, 2990, 2994, 2996, 3004, 3010, 3014, 3016, 3024, 3028: oled_data = 16'b1101110111111110;
    2988, 3006, 3012, 3018, 3022, 3026: oled_data = 16'b1101110110111110;
    2999, 3001, 3029, 3518, 3577, 3585, 3591, 3592, 3668, 3669: oled_data = 16'b1101110111111101;
    3670, 3682, 3971, 4130: oled_data = 16'b1101110111111101;
    3002, 3030: oled_data = 16'b1110010110111110;
    3033, 3076, 3132, 3171, 3229, 3362, 4226, 4419, 4477, 4516: oled_data = 16'b1110011000111101;
    4572, 4616, 4627, 4629, 4633, 4635, 4637, 4639, 4650, 4652: oled_data = 16'b1110011000111101;
    4660, 4663, 4665: oled_data = 16'b1110011000111101;
    3046: oled_data = 16'b1100101110001000;
    3047: oled_data = 16'b1101010000001011;
    3048: oled_data = 16'b1101010010101110;
    3051, 3058, 3148: oled_data = 16'b1110010110110011;
    3052: oled_data = 16'b1101110001001100;
    3053: oled_data = 16'b1101110010101101;
    3054, 3240: oled_data = 16'b1101110100110000;
    3055, 3146, 3152, 3247, 3249, 4015, 4112, 4301, 4396, 4398: oled_data = 16'b1111111101111100;
    4401, 4689, 4780, 4785: oled_data = 16'b1111111101111100;
    3056, 3720: oled_data = 16'b1110111100111010;
    3057, 3536, 3538, 3920, 4109: oled_data = 16'b1110111100111011;
    3059: oled_data = 16'b1101010000001100;
    3060: oled_data = 16'b1101010001001100;
    3061, 3239, 4583: oled_data = 16'b1100101111001010;
    3065: oled_data = 16'b1011101100000101;
    3066: oled_data = 16'b1000101000000100;
    3067: oled_data = 16'b0111001011001010;
    3077, 3131, 3480, 3487, 3554, 3572, 3581, 3650, 3681, 3746: oled_data = 16'b1101110110111101;
    3842, 3938, 4034, 4323, 4381, 4476, 4517, 4571: oled_data = 16'b1101110110111101;
    3078, 3486: oled_data = 16'b1100110010111011;
    3079, 3173: oled_data = 16'b1011001101011001;
    3080, 3094, 3101, 3107, 3116, 3126, 3127: oled_data = 16'b1010001100011000;
    3081, 3087, 3089, 3092, 3093, 3095, 3096, 3100, 3102, 3105: oled_data = 16'b1010101011011000;
    3106, 3109, 3110, 3112, 3115, 3117, 3124, 3125, 4053: oled_data = 16'b1010101011011000;
    3082, 3084, 3086, 3088, 3090, 3098, 3104, 3113, 3119, 3123: oled_data = 16'b1010001011011000;
    4051, 4052, 4054, 4228: oled_data = 16'b1010001011011000;
    3083, 3085, 3091, 3097, 3099, 3103, 3108, 3111, 3114, 3118: oled_data = 16'b1010101100011000;
    3120, 3122, 3128: oled_data = 16'b1010101100011000;
    3121: oled_data = 16'b1010001011011001;
    3129: oled_data = 16'b1010101101011001;
    3130, 3866: oled_data = 16'b1100110010111100;
    3141: oled_data = 16'b1100010011101110;
    3142, 5356: oled_data = 16'b1101110011101100;
    3143: oled_data = 16'b1100001111001010;
    3145, 3154, 3241, 3433, 3439, 3441, 3534, 4881: oled_data = 16'b1111011101111011;
    3149, 4009: oled_data = 16'b1110010100110000;
    3150, 3440: oled_data = 16'b1111011100111011;
    3155, 3437: oled_data = 16'b1111011100111010;
    3156: oled_data = 16'b1101110110110011;
    3158, 4220: oled_data = 16'b1111010100101001;
    3159, 5741: oled_data = 16'b1111011000110000;
    3160, 4390: oled_data = 16'b1111011000110011;
    3162: oled_data = 16'b1010001100000011;
    3163: oled_data = 16'b0111101100001010;
    3172, 3228, 3363, 3974, 4518, 4570: oled_data = 16'b1101010100111101;
    3174, 3269, 3417, 4138: oled_data = 16'b0111000011010011;
    3175, 3225, 3365: oled_data = 16'b0111100101010011;
    3176, 3180, 3186, 3188, 3190, 3191, 3193, 3194, 3196, 3199: oled_data = 16'b1000101000010100;
    3200, 3202, 3203, 3205, 3209, 3211, 3215, 3217, 3219, 3224: oled_data = 16'b1000101000010100;
    3177, 3179, 3181, 3183, 3218, 3220, 3223, 3653, 3845, 4037: oled_data = 16'b1000000111010100;
    3178, 3182, 3184, 3185, 3187, 3189, 3192, 3195, 3198, 3207: oled_data = 16'b1000001000010100;
    3213, 3216, 3221, 3941: oled_data = 16'b1000001000010100;
    3197, 3208, 3212, 3214: oled_data = 16'b1000101000010101;
    3201, 3204, 3206, 3210: oled_data = 16'b1000001000010101;
    3222: oled_data = 16'b1000100111010100;
    3226, 3419: oled_data = 16'b0111000100010011;
    3227, 3275, 3279, 3280, 3282, 3966: oled_data = 16'b1011101110011010;
    3236: oled_data = 16'b0111101100001011;
    3237, 3334, 4582: oled_data = 16'b1011001111001010;
    3238: oled_data = 16'b1101110010101100;
    3244: oled_data = 16'b1110011000110110;
    3245: oled_data = 16'b1101010110110011;
    3246, 4300, 4779: oled_data = 16'b1111111111111101;
    3251: oled_data = 16'b1110111001110101;
    3252: oled_data = 16'b1100110000001100;
    3253: oled_data = 16'b1100101111001001;
    3254: oled_data = 16'b1100001110000111;
    3255, 3740, 4219: oled_data = 16'b1011001100000110;
    3256: oled_data = 16'b1110110111110001;
    3257, 5354: oled_data = 16'b1110010101101101;
    3258: oled_data = 16'b1001001001000011;
    3268, 3324, 3870, 3962, 4475, 4542, 4548, 4559, 4566, 4568: oled_data = 16'b1100010000011011;
    3270: oled_data = 16'b1001001011010101;
    3271, 3366, 3678, 3882, 4569: oled_data = 16'b1100010001011011;
    3272, 3273, 3274, 3276, 3278, 3281, 3285: oled_data = 16'b1011101110011011;
    3277, 3676: oled_data = 16'b1011101101011010;
    3283, 4523, 4525, 4527, 4531, 4533, 4537, 4543, 4545, 4550: oled_data = 16'b1011101111011011;
    4554, 4556, 4560, 4564: oled_data = 16'b1011101111011011;
    3284, 3286, 3287, 3288, 3290, 3291, 3858, 4090, 4186, 4534: oled_data = 16'b1011101111011010;
    4536, 4541, 4547, 4558: oled_data = 16'b1011101111011010;
    3289, 3292, 3294, 3296, 3994: oled_data = 16'b1011001111011010;
    3293, 3295, 3300: oled_data = 16'b1011101111011001;
    3297, 3298, 3299, 3301, 3302, 3303, 3304, 3306, 3307, 3706: oled_data = 16'b1011001111011001;
    3305, 3309, 3610, 3802: oled_data = 16'b1011001111011000;
    3308, 3311, 3514: oled_data = 16'b1010101111011000;
    3310, 3312, 3313, 3314, 3942, 4038: oled_data = 16'b1010101110011000;
    3315, 3317: oled_data = 16'b1010101110010111;
    3316: oled_data = 16'b1010001101011000;
    3318: oled_data = 16'b1010001110011000;
    3319: oled_data = 16'b1010101101010111;
    3320: oled_data = 16'b1010001101010111;
    3321, 4344, 4346, 4349, 4350, 4354: oled_data = 16'b1011010001011001;
    3322: oled_data = 16'b1001001010010101;
    3323: oled_data = 16'b0111000011010010;
    3332, 4415: oled_data = 16'b1011010100110100;
    3333, 5647: oled_data = 16'b1000001011001001;
    3335, 4295, 4391, 4485: oled_data = 16'b1111010111110010;
    3336: oled_data = 16'b1110011000110101;
    3337, 3442, 4207, 4492, 5750: oled_data = 16'b1111011101111100;
    3339, 3435, 3819, 5652: oled_data = 16'b1110011001110111;
    3340, 4022, 4490, 5642: oled_data = 16'b1101111001110111;
    3341: oled_data = 16'b1110011001111000;
    3342, 4214: oled_data = 16'b1101111000110110;
    3347: oled_data = 16'b1110111010111001;
    3349: oled_data = 16'b1110110011101010;
    3351, 5361: oled_data = 16'b1101010011101100;
    3352: oled_data = 16'b1101010010101100;
    3353: oled_data = 16'b1001101011000110;
    3354, 3646, 4125, 4987, 5359, 5455: oled_data = 16'b1000001011001000;
    3361, 3475, 3570, 3588, 3590, 3593, 3597, 4668, 4711: oled_data = 16'b1110111100111110;
    3364, 3601: oled_data = 16'b1001101001010111;
    3367, 3369, 3370, 3372, 3373, 3375, 3376, 3468, 4271, 4272: oled_data = 16'b1001000010011000;
    4273, 4274, 4278, 4280: oled_data = 16'b1001000010011000;
    3368, 3371: oled_data = 16'b1001000001011000;
    3374: oled_data = 16'b1000100001011000;
    3377, 3466, 3467, 3469, 3470, 3566, 3567, 3984, 4080, 4081: oled_data = 16'b1001000011011000;
    4082, 4170, 4178, 4179, 4180, 4181, 4182, 4183: oled_data = 16'b1001000011011000;
    3378, 3568, 3664, 4166, 4168, 4169, 4171, 4175: oled_data = 16'b1001000100011000;
    3379, 3385, 3673, 3677, 3769, 3773, 3970, 4072, 4077: oled_data = 16'b1010000111011001;
    3380, 3382, 3665, 3983, 4067: oled_data = 16'b1010001000011001;
    3381, 3387: oled_data = 16'b1010001000011000;
    3383, 3384, 3389, 3788: oled_data = 16'b1001100111011000;
    3386, 3388, 3393, 4055: oled_data = 16'b1001101000011000;
    3390, 3792, 3961, 4060, 4061, 4167: oled_data = 16'b1001000101010111;
    3391, 3857: oled_data = 16'b1001000110010111;
    3392, 3394, 3398, 3516, 3612, 3708, 3900, 3996, 4092, 4188: oled_data = 16'b1001101000010111;
    3395, 3397, 3692, 3953, 4058: oled_data = 16'b1001100111010111;
    3396: oled_data = 16'b1000100110010111;
    3399: oled_data = 16'b1001101000010110;
    3400: oled_data = 16'b1001001000010111;
    3401, 3404, 3407, 3460, 3652, 3844, 4036, 4132: oled_data = 16'b1001000111010110;
    3402: oled_data = 16'b1000100110010110;
    3403, 3408, 4474: oled_data = 16'b1000100110010101;
    3405, 3406: oled_data = 16'b1001001000010110;
    3409, 3506, 3507, 3509, 3608, 3944, 4141, 4144, 4146, 4243: oled_data = 16'b0111100011010100;
    4244, 4246: oled_data = 16'b0111100011010100;
    3410, 3512, 4136, 4235, 4237, 4238, 4239, 4240: oled_data = 16'b0111000010010011;
    3411, 3412, 3513, 3609, 4039, 4234, 4236: oled_data = 16'b0111000001010011;
    3414: oled_data = 16'b0111000001010010;
    3418, 4334, 4335, 4337: oled_data = 16'b1011010000011000;
    3420, 3695: oled_data = 16'b1010001010011000;
    3427: oled_data = 16'b1010101101001100;
    3428: oled_data = 16'b1100101110001101;
    3429, 5544: oled_data = 16'b1000001011001010;
    3430: oled_data = 16'b1001010001001111;
    3431, 3628: oled_data = 16'b1101110110110000;
    3436: oled_data = 16'b1110011010111000;
    3438: oled_data = 16'b1101010111110101;
    3443, 4586, 4682: oled_data = 16'b1111011011111000;
    3444: oled_data = 16'b1111011001110001;
    3447: oled_data = 16'b1110010101101111;
    3448: oled_data = 16'b1001101011000101;
    3449, 5263: oled_data = 16'b0111101010001000;
    3459, 3517, 4131: oled_data = 16'b1101010011111101;
    3461, 3749, 4133: oled_data = 16'b1000001000010011;
    3462: oled_data = 16'b1011001101011010;
    3463, 3561, 3562, 3659, 3660, 3662, 3988, 3990, 4087, 4263: oled_data = 16'b1000100010010111;
    3464, 3564, 3985, 4184, 4267, 4269: oled_data = 16'b1001000011010111;
    3465, 4084: oled_data = 16'b1000100011011000;
    3471: oled_data = 16'b1001100011011001;
    3472, 4076: oled_data = 16'b1001100100011001;
    3473, 3869, 4071: oled_data = 16'b1001100110011001;
    3474: oled_data = 16'b1100110000011011;
    3491, 3954: oled_data = 16'b1110111011111101;
    3492: oled_data = 16'b1100110011111011;
    3493, 3584, 3680, 4614: oled_data = 16'b1110011001111101;
    3498: oled_data = 16'b1100110100111011;
    3499, 3688: oled_data = 16'b1101110110111100;
    3505: oled_data = 16'b1010001100010111;
    3508, 3604, 3605, 3606, 3607, 3703, 3945, 4040, 4042, 4043: oled_data = 16'b0111100010010100;
    4044, 4045, 4046, 4142, 4143, 4241, 4242, 4249: oled_data = 16'b0111100010010100;
    3510: oled_data = 16'b0111000010010100;
    3511: oled_data = 16'b0111100011010011;
    3515, 3557, 3803: oled_data = 16'b1000000111010011;
    3521: oled_data = 16'b1100011001111001;
    3522: oled_data = 16'b1010001011001010;
    3523: oled_data = 16'b1111010000001110;
    3524: oled_data = 16'b1110101110001101;
    3525: oled_data = 16'b1100001000000111;
    3526: oled_data = 16'b1001000110000101;
    3527, 5743: oled_data = 16'b0111101010000111;
    3529: oled_data = 16'b1101010111110100;
    3530, 3722, 5745: oled_data = 16'b1100110111110110;
    3531, 4118, 4406: oled_data = 16'b1101111000110101;
    3532: oled_data = 16'b1110111011110111;
    3533, 4028: oled_data = 16'b1110111011111010;
    3540: oled_data = 16'b1111010011100110;
    3542: oled_data = 16'b1101010110110000;
    3545, 4222: oled_data = 16'b1011110101110101;
    3549, 3643, 4031, 5448: oled_data = 16'b1110011011111010;
    3555, 3709, 3843, 4035: oled_data = 16'b1101010010111101;
    3556, 3804: oled_data = 16'b1001000111010111;
    3558: oled_data = 16'b1011001110011010;
    3559: oled_data = 16'b1000100001010110;
    3560, 3563, 3661, 3759, 3890, 3986, 3987, 3989, 4086, 4088: oled_data = 16'b1000100011010111;
    4159, 4261, 4262, 4264, 4266: oled_data = 16'b1000100011010111;
    3565, 4268, 4270: oled_data = 16'b1000100010011000;
    3569: oled_data = 16'b1010101000011001;
    3575: oled_data = 16'b1101010101111101;
    3582, 3595, 3600, 3693, 3789, 3861: oled_data = 16'b1101010101111100;
    3599: oled_data = 16'b1101111000111100;
    3602, 3603, 3698, 3699, 3701, 3796, 3800, 3848, 3850, 3949: oled_data = 16'b1000000011010101;
    3951, 4048, 4145, 4245, 4251: oled_data = 16'b1000000011010101;
    3615: oled_data = 16'b1100110111111011;
    3616: oled_data = 16'b1010101110001110;
    3617: oled_data = 16'b1001101000001000;
    3618: oled_data = 16'b1011101010001001;
    3619: oled_data = 16'b1110110111110100;
    3620: oled_data = 16'b1110010000001111;
    3621: oled_data = 16'b1010000010000000;
    3622: oled_data = 16'b1010000110000001;
    3623: oled_data = 16'b1001001110001010;
    3624: oled_data = 16'b1010010101110101;
    3626, 4506: oled_data = 16'b0110101001001000;
    3627: oled_data = 16'b1011001110000101;
    3633, 4017, 4099, 5271, 5746: oled_data = 16'b1110011100111100;
    3635, 3731, 3932, 4018, 4124: oled_data = 16'b1110111000110010;
    3636: oled_data = 16'b1101010000000011;
    3638, 3735: oled_data = 16'b0110101001000110;
    3639: oled_data = 16'b0111001001000111;
    3644, 3645: oled_data = 16'b1000101100001001;
    3647, 4319: oled_data = 16'b1011110100110011;
    3655, 3752, 3753, 3795, 3853, 3893, 3895, 3993, 4253, 4256: oled_data = 16'b1000000010010110;
    4257, 4259: oled_data = 16'b1000000010010110;
    3656, 3657, 3794, 3855, 3892, 3991, 4156, 4158, 4160, 4260: oled_data = 16'b1000100011010110;
    3658, 3756, 3758, 3891, 3992, 4258: oled_data = 16'b1000100010010110;
    3663, 3889, 4057, 4161, 4162: oled_data = 16'b1000100100010111;
    3671, 3901, 4324, 4380: oled_data = 16'b1100110001011100;
    3672, 3979, 4078: oled_data = 16'b1010101001011010;
    3674, 3770: oled_data = 16'b1101010011111100;
    3691: oled_data = 16'b1010101100011001;
    3696: oled_data = 16'b1000100101010110;
    3697, 3793, 3856, 4149, 4151, 4153, 4157: oled_data = 16'b1000100100010110;
    3700, 3702, 3946, 4248, 4252: oled_data = 16'b0111100010010101;
    3704, 3947, 4047: oled_data = 16'b0111100011010101;
    3705, 3847, 3943: oled_data = 16'b0111100001010100;
    3707, 4091: oled_data = 16'b0111100110010011;
    3710: oled_data = 16'b1100110110111100;
    3711: oled_data = 16'b1000101000001000;
    3712: oled_data = 16'b1100100010000000;
    3713: oled_data = 16'b1101100010000001;
    3714, 3809: oled_data = 16'b1101000011000010;
    3715: oled_data = 16'b0111101101000100;
    3716: oled_data = 16'b1001000111000100;
    3717: oled_data = 16'b1101001011001010;
    3718: oled_data = 16'b1101001100001001;
    3719: oled_data = 16'b1011101000000100;
    3721, 5732, 5733, 5753: oled_data = 16'b1011010110110110;
    3723: oled_data = 16'b1110011100111010;
    3724, 3817, 4013, 5176, 5256, 5352: oled_data = 16'b1110111100111100;
    3726, 5663, 5739, 5924: oled_data = 16'b1101111011111011;
    3734, 4504: oled_data = 16'b1101110010101000;
    3739, 4892: oled_data = 16'b1000101011001001;
    3741, 4508: oled_data = 16'b1110010011101001;
    3743: oled_data = 16'b1010101111001000;
    3747, 3997: oled_data = 16'b1100110010111101;
    3748, 3940: oled_data = 16'b1001000110010110;
    3751, 3801: oled_data = 16'b0111100001010101;
    3754, 3755, 3757, 3854, 3894, 3896, 3952, 4154, 4155, 4255: oled_data = 16'b1000000011010110;
    3760, 3888, 3965, 4163, 4164, 4165: oled_data = 16'b1001000100010111;
    3761, 3865, 3884, 3969, 4064: oled_data = 16'b1001100110011000;
    3762: oled_data = 16'b1100010010111011;
    3768, 3864, 3868, 3968: oled_data = 16'b1011001100011010;
    3772: oled_data = 16'b1011001100011011;
    3774: oled_data = 16'b1100110000011100;
    3786, 3859, 3879, 3976: oled_data = 16'b1101010100111100;
    3787: oled_data = 16'b1010001001011001;
    3791: oled_data = 16'b1010101010011000;
    3797, 3798, 3799, 3849, 3851, 3852, 3897, 3948, 3950, 4247: oled_data = 16'b1000000010010101;
    4250, 4254: oled_data = 16'b1000000010010101;
    3805: oled_data = 16'b1101110011111110;
    3806: oled_data = 16'b1010010001010110;
    3807: oled_data = 16'b1010000100000011;
    3808: oled_data = 16'b1110000011000010;
    3810: oled_data = 16'b1101100100000010;
    3811: oled_data = 16'b1001000111000010;
    3812, 4699: oled_data = 16'b1001101101000111;
    3813: oled_data = 16'b1110101111001110;
    3814: oled_data = 16'b1110110001001111;
    3815: oled_data = 16'b1101101011001011;
    3816: oled_data = 16'b1110111011111011;
    3818: oled_data = 16'b1011001110001010;
    3826, 4486: oled_data = 16'b1111111010110101;
    3828, 4311, 4407, 5357: oled_data = 16'b1111010110101100;
    3829: oled_data = 16'b1101111000110011;
    3831: oled_data = 16'b1011001100000101;
    3832: oled_data = 16'b1001001011001000;
    3833, 5832, 5834, 5844, 5846: oled_data = 16'b1100111000110111;
    3834, 4967, 5946: oled_data = 16'b1101011001111001;
    3835: oled_data = 16'b0110101001000101;
    3846: oled_data = 16'b1010101110011001;
    3860: oled_data = 16'b1101010110111100;
    3862: oled_data = 16'b1110111001111101;
    3872: oled_data = 16'b1100010000011100;
    3874: oled_data = 16'b1011101100011011;
    3883, 3964, 4070: oled_data = 16'b1010101001011001;
    3885: oled_data = 16'b1101110101111100;
    3887: oled_data = 16'b1010001010011001;
    3899, 4187: oled_data = 16'b0111100111010011;
    3902: oled_data = 16'b1001110010110100;
    3903: oled_data = 16'b1100110011110010;
    3904: oled_data = 16'b1101000101000100;
    3905: oled_data = 16'b1101100011000010;
    3906: oled_data = 16'b1101000011000001;
    3907: oled_data = 16'b1110101110001111;
    3908, 4005: oled_data = 16'b1110111000111000;
    3909: oled_data = 16'b1101101010001001;
    3910: oled_data = 16'b1110001100001011;
    3911: oled_data = 16'b1101110011110010;
    3914: oled_data = 16'b1010001100000110;
    3915, 4890: oled_data = 16'b1110111000110100;
    3923: oled_data = 16'b1111110101100111;
    3924, 4694, 4792, 5068: oled_data = 16'b1111010111101111;
    3925: oled_data = 16'b1101111010111000;
    3926: oled_data = 16'b1110011000110001;
    3927: oled_data = 16'b1101110001001001;
    3928: oled_data = 16'b0111101010000101;
    3929: oled_data = 16'b1000001101001101;
    3930: oled_data = 16'b1010110001001110;
    3931, 4409: oled_data = 16'b1001101011000111;
    3933: oled_data = 16'b1011110001001010;
    3934: oled_data = 16'b1010001111001100;
    3935, 4511: oled_data = 16'b1010110011110001;
    3959: oled_data = 16'b1110111010111101;
    3960, 4059, 4063: oled_data = 16'b1010001001011000;
    3975: oled_data = 16'b1010101000011010;
    3980, 4066: oled_data = 16'b1001100101011000;
    3981: oled_data = 16'b1100110011111100;
    3998: oled_data = 16'b1011110011110101;
    4000, 5064: oled_data = 16'b1101010111110111;
    4001: oled_data = 16'b1101010010110001;
    4002: oled_data = 16'b1101010101110101;
    4003, 4014, 5160, 5738, 5748: oled_data = 16'b1110111101111100;
    4006: oled_data = 16'b1110110111110111;
    4010, 4384: oled_data = 16'b1101010010101001;
    4011, 4210, 4509: oled_data = 16'b1111011010110100;
    4012: oled_data = 16'b1110011101111101;
    4020, 4503: oled_data = 16'b1110010100101001;
    4021: oled_data = 16'b1101110110101111;
    4023: oled_data = 16'b1110110110101100;
    4024, 4213: oled_data = 16'b1010101100000110;
    4025: oled_data = 16'b0110100111000101;
    4026: oled_data = 16'b1000001010000101;
    4027: oled_data = 16'b1110010100101011;
    4030: oled_data = 16'b1001101111001110;
    4041, 4140: oled_data = 16'b0111000011010100;
    4050: oled_data = 16'b1001101001011000;
    4056: oled_data = 16'b1000100101010111;
    4062: oled_data = 16'b1001000110011000;
    4065: oled_data = 16'b1001000101011000;
    4068: oled_data = 16'b1010101010011001;
    4069, 4073, 4074: oled_data = 16'b1010101010011010;
    4075: oled_data = 16'b1010000110011001;
    4079: oled_data = 16'b1001100101011001;
    4083, 4085, 4265: oled_data = 16'b1001000010010111;
    4089, 4185: oled_data = 16'b1000100001010111;
    4093: oled_data = 16'b1101110011111111;
    4094: oled_data = 16'b1010010000010010;
    4095: oled_data = 16'b1011110000001001;
    4096, 5837: oled_data = 16'b1101011000110110;
    4097, 5937, 5941, 5949: oled_data = 16'b1100111010111001;
    4098: oled_data = 16'b1101011011111001;
    4103: oled_data = 16'b1111011001110111;
    4104, 4296: oled_data = 16'b1110110101110000;
    4105: oled_data = 16'b1111010110110001;
    4106, 4195: oled_data = 16'b1100110001001011;
    4107: oled_data = 16'b1110111010110101;
    4115, 4308: oled_data = 16'b1110110010100101;
    4116: oled_data = 16'b1100001111000011;
    4119, 4692: oled_data = 16'b1110110101101011;
    4122: oled_data = 16'b1000101011000111;
    4126, 4575, 4989, 5084, 5842: oled_data = 16'b1100111000111000;
    4134: oled_data = 16'b1010101101011000;
    4147, 4148, 4150: oled_data = 16'b1000000100010101;
    4172: oled_data = 16'b1001100100011000;
    4173: oled_data = 16'b1001000100011001;
    4174, 4176: oled_data = 16'b1001100011011000;
    4177: oled_data = 16'b1001000011011001;
    4189: oled_data = 16'b1101010100111110;
    4190: oled_data = 16'b1100010011110111;
    4191, 4480: oled_data = 16'b1100010000000111;
    4192: oled_data = 16'b1100110001001001;
    4193, 4196: oled_data = 16'b1100110011101101;
    4194: oled_data = 16'b1100110011101110;
    4198: oled_data = 16'b1110110011101111;
    4199: oled_data = 16'b1110110011101110;
    4201: oled_data = 16'b1111010101110000;
    4202: oled_data = 16'b1100010010101101;
    4203: oled_data = 16'b1110111010110110;
    4211, 4216, 4600, 4969, 5077: oled_data = 16'b1110110100101000;
    4215: oled_data = 16'b1110010101101011;
    4217, 4601: oled_data = 16'b1011010000001001;
    4218, 4698: oled_data = 16'b1000001010000111;
    4221: oled_data = 16'b1000001101001001;
    4227: oled_data = 16'b1101110100111101;
    4229: oled_data = 16'b0110100100010010;
    4230, 4328, 4332, 4336, 4338, 4339, 4341, 4342, 4343, 4345: oled_data = 16'b1011010001011000;
    4231: oled_data = 16'b1000000101010100;
    4232: oled_data = 16'b0110100010010010;
    4233: oled_data = 16'b0110100010010011;
    4275, 4276, 4279: oled_data = 16'b1001000010011001;
    4277: oled_data = 16'b1001100010011000;
    4281: oled_data = 16'b1010000111011010;
    4282, 4352, 4353, 4355, 4357, 4358, 4359, 4360, 4361, 4365: oled_data = 16'b1011110001011001;
    4367: oled_data = 16'b1011110001011001;
    4283: oled_data = 16'b0110100011010001;
    4284: oled_data = 16'b1010101011011001;
    4286: oled_data = 16'b1101010111111100;
    4288, 4289, 4386, 4604: oled_data = 16'b1100110000000111;
    4290: oled_data = 16'b1100110001001000;
    4292: oled_data = 16'b1101110001001010;
    4293: oled_data = 16'b1110110100101110;
    4294: oled_data = 16'b1110110100101111;
    4297: oled_data = 16'b1111110111110001;
    4298: oled_data = 16'b1101010101110001;
    4299: oled_data = 16'b1110011010111001;
    4307: oled_data = 16'b1110010111110001;
    4310: oled_data = 16'b1101111001110101;
    4314, 4602, 4893, 5366, 5558: oled_data = 16'b0110101001000111;
    4317: oled_data = 16'b1111011011110110;
    4318: oled_data = 16'b1001101111001101;
    4325: oled_data = 16'b0111100100010011;
    4326, 4430: oled_data = 16'b0111100111010010;
    4327: oled_data = 16'b1011010010111000;
    4329, 4331: oled_data = 16'b1011010000010111;
    4330: oled_data = 16'b1010110001011000;
    4333: oled_data = 16'b1010110000011000;
    4340, 4347: oled_data = 16'b1011010000011001;
    4348: oled_data = 16'b1011110001011000;
    4351, 4356, 4363: oled_data = 16'b1011110000011001;
    4362, 4364, 4366, 4368, 4369, 4371, 4373, 4375: oled_data = 16'b1011110001011010;
    4370, 4372, 4374, 4376: oled_data = 16'b1100010001011010;
    4377: oled_data = 16'b1011110010111001;
    4378, 4448, 4454, 4458, 4461, 4466, 4469: oled_data = 16'b0111000110010001;
    4382: oled_data = 16'b1101111001111101;
    4383: oled_data = 16'b1010110000001100;
    4385, 4697: oled_data = 16'b1100001111000111;
    4387: oled_data = 16'b1100110001001010;
    4392, 4403, 4787: oled_data = 16'b1111111001110011;
    4393: oled_data = 16'b1101010011101111;
    4394: oled_data = 16'b1010010001001110;
    4404: oled_data = 16'b1110110011100101;
    4405: oled_data = 16'b1101010010100111;
    4408: oled_data = 16'b1101110000000110;
    4411: oled_data = 16'b0110101000000101;
    4414, 4984: oled_data = 16'b1010001110001000;
    4421, 4520, 4529, 4562: oled_data = 16'b1011110000011011;
    4422: oled_data = 16'b1000000110010100;
    4423, 4473: oled_data = 16'b0110100100010001;
    4424, 4425, 4427, 4429, 4432, 4434, 4435, 4437, 4438, 4440: oled_data = 16'b0111100110010010;
    4441, 4444, 4450, 4459, 4462: oled_data = 16'b0111100110010010;
    4426, 4428, 4431, 4433, 4436, 4439, 4443, 4445, 4447, 4449: oled_data = 16'b0111000110010010;
    4451, 4452, 4453, 4455, 4456, 4457, 4460, 4463, 4465, 4468: oled_data = 16'b0111000110010010;
    4470, 4471, 4472: oled_data = 16'b0111000110010010;
    4442, 4446, 4464, 4467: oled_data = 16'b0111100110010001;
    4479: oled_data = 16'b1011110011110000;
    4481, 4484: oled_data = 16'b1101110100101100;
    4482: oled_data = 16'b1101010011101011;
    4483: oled_data = 16'b1101010011101010;
    4487: oled_data = 16'b1111111001110100;
    4488: oled_data = 16'b1100110001001101;
    4489: oled_data = 16'b0111100111000100;
    4500: oled_data = 16'b1110110101101010;
    4501: oled_data = 16'b1101110110110001;
    4502: oled_data = 16'b1101110101101101;
    4505: oled_data = 16'b1011001110001000;
    4507: oled_data = 16'b0111001001000110;
    4519: oled_data = 16'b1100110001011011;
    4521, 4535, 4538, 4540, 4551, 4553, 4557, 4563: oled_data = 16'b1100001111011011;
    4522, 4539: oled_data = 16'b1011110000011010;
    4524, 4532, 4555: oled_data = 16'b1100010000011010;
    4526, 4528, 4530, 4544, 4546, 4549, 4552, 4561, 4565, 4567: oled_data = 16'b1100001111011010;
    4576: oled_data = 16'b1000101110001011;
    4578: oled_data = 16'b1011001111001000;
    4584: oled_data = 16'b1010101100000101;
    4585: oled_data = 16'b1101010001001000;
    4589, 4686, 4783, 4875, 4877, 4880: oled_data = 16'b1111111101111101;
    4597: oled_data = 16'b1101111001110110;
    4603: oled_data = 16'b0110101000000110;
    4605: oled_data = 16'b1111010111110000;
    4607: oled_data = 16'b1010110011110011;
    4612: oled_data = 16'b1111011011111111;
    4648: oled_data = 16'b1101111000111101;
    4662: oled_data = 16'b1101111000111110;
    4673, 5636, 5731, 5925, 5928, 5930, 5931, 5932, 5933, 5938: oled_data = 16'b1100111001111001;
    5939, 5940, 5942, 5945, 5947, 5950: oled_data = 16'b1100111001111001;
    4674: oled_data = 16'b1010010010110001;
    4675: oled_data = 16'b1011010011110000;
    4677: oled_data = 16'b1010001101000111;
    4678: oled_data = 16'b1010001101000110;
    4679: oled_data = 16'b1010101101001001;
    4680: oled_data = 16'b1011101111000101;
    4693: oled_data = 16'b1101111010110111;
    4701, 5072: oled_data = 16'b1111110111101110;
    4703, 5638: oled_data = 16'b1010110011110010;
    4773: oled_data = 16'b1011110101110100;
    4776: oled_data = 16'b0110001000000110;
    4778, 5451: oled_data = 16'b1110111010111000;
    4788: oled_data = 16'b1111010110101011;
    4789: oled_data = 16'b1110011000110100;
    4790: oled_data = 16'b1101111000110100;
    4791, 4797: oled_data = 16'b1101011000110100;
    4793: oled_data = 16'b1101110011101011;
    4794: oled_data = 16'b1101010000001001;
    4874: oled_data = 16'b1111011100110111;
    4889, 5740: oled_data = 16'b1110011011111001;
    4891: oled_data = 16'b1101110011101001;
    4981, 4983, 5078, 5172: oled_data = 16'b1101110001000101;
    4982: oled_data = 16'b1101010001000100;
    4985, 5735: oled_data = 16'b1000001101001011;
    4988, 5545: oled_data = 16'b0110001001000110;
    5075: oled_data = 16'b1110110100100111;
    5079: oled_data = 16'b1001001011000101;
    5080: oled_data = 16'b1011110100110010;
    5082: oled_data = 16'b1101011000111000;
    5167: oled_data = 16'b1011110000001000;
    5168: oled_data = 16'b1011110000000111;
    5171: oled_data = 16'b1101110010100110;
    5174: oled_data = 16'b1011001111000111;
    5175: oled_data = 16'b1011010011110001;
    5257: oled_data = 16'b1000101101001010;
    5258: oled_data = 16'b1100110000000110;
    5260: oled_data = 16'b1101010000000101;
    5262: oled_data = 16'b1100010000000101;
    5264: oled_data = 16'b0110001000001000;
    5265: oled_data = 16'b1100010000000110;
    5266: oled_data = 16'b1101010000000100;
    5267: oled_data = 16'b1100001101000100;
    5268, 5742: oled_data = 16'b1100101111000100;
    5269: oled_data = 16'b1100001111000101;
    5270: oled_data = 16'b0111001010001000;
    5355: oled_data = 16'b1101010010101011;
    5360, 5648: oled_data = 16'b0101100111000110;
    5362: oled_data = 16'b1110010100101100;
    5363: oled_data = 16'b1011101110001011;
    5365: oled_data = 16'b1100110000000100;
    5450: oled_data = 16'b1100110110110100;
    5453: oled_data = 16'b1110011000110010;
    5456: oled_data = 16'b0101100111000101;
    5457: oled_data = 16'b1011110101110010;
    5459: oled_data = 16'b1110011011111000;
    5462, 5551: oled_data = 16'b0111101011001000;
    5546: oled_data = 16'b1010101100000111;
    5548: oled_data = 16'b1101010001001001;
    5552: oled_data = 16'b0101101000000110;
    5553: oled_data = 16'b1001001010000110;
    5555: oled_data = 16'b1101110010101010;
    5559: oled_data = 16'b1101111010111011;
    5637: oled_data = 16'b1011111000111000;
    5639: oled_data = 16'b1010110010110000;
    5641: oled_data = 16'b1011110110110101;
    5643: oled_data = 16'b1101011000110111;
    5644: oled_data = 16'b1110010110101111;
    5649: oled_data = 16'b1100010101110010;
    5650: oled_data = 16'b1110111010110111;
    5651: oled_data = 16'b1110011001110110;
    5653: oled_data = 16'b1101011000110101;
    5654: oled_data = 16'b1101011001110111;
    5656: oled_data = 16'b1010010011110011;
    5657: oled_data = 16'b1100011000111000;
    5658, 5659, 5661, 5662, 5759, 5833, 5835, 5843, 5845, 5855: oled_data = 16'b1011110111110111;
    5744: oled_data = 16'b0101000111000101;
    5749, 5926, 5927, 5935, 5943, 5944: oled_data = 16'b1101011010111010;
    5752, 5831: oled_data = 16'b1000110000001111;
    5754, 5756, 5758, 5829, 5850, 5851, 5852, 5853: oled_data = 16'b1010110101110101;
    5755, 5828, 5849: oled_data = 16'b1010110110110110;
    5757: oled_data = 16'b1010110110110101;
    5830: oled_data = 16'b1001010001010001;
    5836: oled_data = 16'b1100111000111001;
    5838: oled_data = 16'b1011110010101100;
    5840: oled_data = 16'b0111101101001100;
    5847: oled_data = 16'b1000101111001110;
    5848: oled_data = 16'b1001110010110010;
    5854: oled_data = 16'b1010110100110101;
    5929: oled_data = 16'b1100111001111010;
    5934: oled_data = 16'b1100111010111011;
    5936: oled_data = 16'b1101011010111011;
    5948: oled_data = 16'b1101011001111010;
    default: oled_data = 16'b0000000000000000;
    endcase
    end

endmodule
