`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.10.2024 15:23:34
// Design Name: 
// Module Name: frame_data_feature2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// feature 3 - level 1
module frame_data_feature3( 
    input CLOCK,
    output reg [6:0] seg,
    output reg [3:0] an,
    output reg [1:0] lives_level,
    output reg [15:0] oled_data,
    output reg [1:0] level_completed,
    output reg [1:0] level0_completed,
    output reg [1:0] level1_completed,
    output reg [1:0] level2_completed,
    output reg [1:0] tryagain,
    input frame_rate, 
    input [12:0] pixel_index,  
    input [1:0] pointer_clk,
    input [15:0] x_min,
    input fast_clk,
    input [15:0] x_max,
    input [3:0] state,
    input btnC
    );
    
    always @(posedge CLOCK) begin
          if (state == 4'b0011) begin
          if (level1_completed) begin
              // Third level
              seg <= 7'b0110000;  
              an <= 4'b0000;      
          end else if (level0_completed) begin
              // second level
              seg <= 7'b0100100;  
              an <= 4'b0000;      
          end else begin
              // first level
              seg <= 7'b1001111;  
              an <= 4'b0000;     
          end end 
          else begin
            an <= 4'b1111;
            seg <= 7'b1111111;
          end
          end

    // moving direction
    reg [1:0] move_dir = 1; // initialized to move right
    reg [6:0] x_pos = 26; // current x-position of the pointer
    reg [6:0] y_pos = 25; // current y-position of the pointer
    
    initial begin
        lives_level <= 3;
        level0_completed <= 0;
        level1_completed <= 0;
        level2_completed <= 0;
        level_completed <= 0;
        tryagain <= 0;
    end

         
    // for debouncing
    reg [7:0] debounce_btnC = 0;
    reg btnC_pressed = 0;
    reg btnC_prev = 0;
    reg btnC_released = 1;
    
    always @(posedge fast_clk) begin
        if (btnC && !btnC_prev && debounce_btnC == 0 && btnC_released) begin
            btnC_pressed <= 1;
            debounce_btnC <= 200;
            btnC_released <= 0;
        end else if (debounce_btnC > 0) begin
            debounce_btnC <= debounce_btnC - 1;
            btnC_pressed <= 0;
        end else if (!btnC) begin
            btnC_released <= 1;
        end else begin
            btnC_pressed <= 0;
        end
            btnC_prev <= btnC;
    end
     
    wire [7:0] x;
    wire [6:0] y;
    assign x = pixel_index % 96;
    assign y = pixel_index / 96;
      
    always @(posedge pointer_clk) begin
        case(move_dir)
            1: // right
                if (x_pos < 70)
                    x_pos <= x_pos + 1;
            2: // left
                if (x_pos > 25)
                x_pos <= x_pos - 1;
        endcase
    end

    
    always@ (posedge frame_rate) begin
        if (x_pos == 70) begin
            move_dir <= 2;
        end else if (x_pos == 25) begin
            move_dir <= 1;
        end 
    end


    // green part of temp bar
    reg is_within_green_area;
    
    always @(posedge fast_clk) begin
    if (state == 4'b0011) begin
        if ((x_pos >= x_min && x_pos <= x_max) &&
            (y_pos >= 22 && y_pos <= 29)) begin
            is_within_green_area <= 1;
    end else begin
            is_within_green_area <= 0;
    end
    
    if (btnC_pressed && is_within_green_area) begin
        level_completed <= level_completed + 1;
    end if (btnC_pressed && !is_within_green_area) begin
        lives_level <= lives_level - 1;
    end end

      
    if (level_completed == 0) begin
         level0_completed <= 0;
         level1_completed <= 0;
         level2_completed <= 0;
         tryagain <= 0;
    end else if (level_completed == 1) begin
         level0_completed <= 1; // first level
         level1_completed <= 0;
         level2_completed <= 0;
         tryagain <= 0;
    end else if (level_completed == 2) begin
         level1_completed <= 1; // second level
         level0_completed <= 0;
         level2_completed <= 0;
         tryagain <= 0;
    end else if (level_completed == 3) begin
         level1_completed <= 0; // third level
         level0_completed <= 0;
         level2_completed <= 1;
         tryagain <= 0;
    end 

    if (lives_level == 0 && !tryagain) begin
        level_completed <= 0;
        level0_completed <= 0;
        level1_completed <= 0;
        level2_completed <= 0;
        tryagain <= 1; 
    end if (btnC_pressed && tryagain) begin
         lives_level <= 3;
         tryagain <= 0;  
    end end   

    // lives
    always @ (posedge frame_rate) begin
        if (lives_level == 3) begin if 
            ((((x == 3 | x == 4 | x == 6 | x == 7) && y == 2)
            | ((x >= 2 && x <= 8) && (y == 3 | y == 4))
            | ((x >= 3 && x <= 7) && y == 5)
            | ((x >= 4 && x <= 6) && y == 6)
            | (x == 5 && y == 7))
            //2nd heart   
            | (((x == 11 | x == 12 | x == 14 | x == 15) && y == 2)
            | ((x >= 10 && x <= 16) && (y == 3 | y == 4))
            | ((x >= 11 && x <= 15) && y == 5)
            | ((x >= 12 && x <= 14) && y == 6)
            | (x == 13 && y == 7))
            //3rd heart
            | (((x == 19 | x == 20 | x == 22 | x == 23) && y == 2)
            | ((x >= 18 && x <= 24) && (y == 3 | y == 4))
            | ((x >= 19 && x <= 23) && y == 5)
            | ((x >= 20 && x <= 22) && y == 6)
            | (x == 21 && y == 7)))
            begin
                oled_data <= 16'b11100_000000_01001;
            end end else if (lives_level == 2) begin if 
            ((((x == 3 | x == 4 | x == 6 | x == 7) && y == 2)
            | ((x >= 2 && x <= 8) && (y == 3 | y == 4))
            | ((x >= 3 && x <= 7) && y == 5)
            | ((x >= 4 && x <= 6) && y == 6)
            | (x == 5 && y == 7))
            //2nd heart   
            | (((x == 11 | x == 12 | x == 14 | x == 15) && y == 2)
            | ((x >= 10 && x <= 16) && (y == 3 | y == 4))
            | ((x >= 11 && x <= 15) && y == 5)
            | ((x >= 12 && x <= 14) && y == 6)
            | (x == 13 && y == 7))
            //3rd heart
            | (((x == 19 | x == 20 | x == 22 | x == 23) && y == 2)
            | ((x == 18 | x == 21 | x == 24) && y == 3)
            | ((x == 18 | x == 24) && y == 4)
            | ((x == 19 | x == 23) && y == 5)
            | ((x == 20 | x == 22) && y == 6)
            | (x == 21 && y == 7)))
            begin
                oled_data <= 16'b11100_000000_01001;
            end end else if (lives_level == 1) begin if 
            ((((x == 3 | x == 4 | x == 6 | x == 7) && y == 2)
            | ((x >= 2 && x <= 8) && (y == 3 | y == 4))
            | ((x >= 3 && x <= 7) && y == 5)
            | ((x >= 4 && x <= 6) && y == 6)
            | (x == 5 && y == 7))
            //2nd heart   
            | (((x == 11 | x == 12 | x == 14 | x == 15) && y == 2)
            | ((x == 10 | x == 13 | x == 16) && y == 3)
            | ((x == 10 | x == 16) && y == 4)
            | ((x == 11 | x == 15) && y == 5)
            | ((x == 12 | x == 14) && y == 6)
            | (x == 13 && y == 7))
            //3rd heart
            | (((x == 19 | x == 20 | x == 22 | x == 23) && y == 2)
            | ((x == 18 | x == 21 | x == 24) && y == 3)
            | ((x == 18 | x == 24) && y == 4)
            | ((x == 19 | x == 23) && y == 5)
            | ((x == 20 | x == 22) && y == 6)
            | (x == 21 && y == 7)))
            begin
                oled_data <= 16'b11100_000000_01001;
            end end

    // draw out black pointer
    if ((x >= x_pos) && (x <= x_pos + 1) && (y >= 25) && (y <= 29)) begin
        oled_data <= 16'b00000_000000_00000;  // black pointer
    end

    // temperature bar
    // red part is ((x >= 24 && x <= 71) && (y >= 22 && y <= 29))
    else if ((x >= x_min && x <= x_max) && (y >= 22 && y <= 29)) oled_data = 16'b0011110011100111; // green part
    else if ((x >= 24 && x <= 71) && (y >= 22 && y <= 29)) oled_data = 16'b1011100010100011; // red part  
        
// background
    else begin
    case (pixel_index)
         0, 1, 7, 8, 9, 14, 15, 16, 17, 22: oled_data = 16'b1111111000111011;
         23, 24, 31, 32, 33, 38, 39, 40, 47, 48: oled_data = 16'b1111111000111011;
         49, 55, 56, 57, 62, 63, 64, 71, 72, 73: oled_data = 16'b1111111000111011;
         79, 80, 81, 86, 87, 88, 95, 102, 104, 111: oled_data = 16'b1111111000111011;
         119, 128, 135, 136, 143, 152, 159, 160, 161, 168: oled_data = 16'b1111111000111011;
         175, 184, 191, 576, 577, 583, 585, 591, 592, 593: oled_data = 16'b1111111000111011;
         598, 600, 601, 607, 608, 609, 615, 616, 617, 623: oled_data = 16'b1111111000111011;
         625, 631, 632, 639, 641, 647, 649, 655, 656, 657: oled_data = 16'b1111111000111011;
         663, 664, 665, 670, 671, 672, 680, 681, 686, 687: oled_data = 16'b1111111000111011;
         689, 695, 696, 703, 705, 710, 711, 713, 719, 720: oled_data = 16'b1111111000111011;
         721, 727, 729, 735, 736, 743, 744, 751, 752, 759: oled_data = 16'b1111111000111011;
         761, 768, 769, 775, 777, 782, 783, 784, 785, 790: oled_data = 16'b1111111000111011;
         791, 792, 799, 800, 808, 809, 815, 817, 823, 824: oled_data = 16'b1111111000111011;
         825, 830, 831, 832, 833, 840, 846, 848, 849, 854: oled_data = 16'b1111111000111011;
         855, 856, 863, 864, 871, 872, 896, 903, 911, 912: oled_data = 16'b1111111000111011;
         919, 921, 927, 929, 936, 943, 944, 952, 958, 959: oled_data = 16'b1111111000111011;
         1344, 1351, 1352, 1353, 1358, 1360, 1367, 1368, 1375, 1377: oled_data = 16'b1111111000111011;
         1382, 1384, 1391, 1393, 1399, 1400, 1407, 1409, 1415, 1416: oled_data = 16'b1111111000111011;
         1423, 1424, 1425, 1431, 1432, 1439, 1440, 1441, 1446, 1448: oled_data = 16'b1111111000111011;
         1454, 1456, 1457, 1462, 1464, 1465, 1471, 1472, 1473, 1479: oled_data = 16'b1111111000111011;
         1481, 1487, 1488, 1494, 1495, 1496, 1497, 1502, 1504, 1505: oled_data = 16'b1111111000111011;
         1511, 1513, 1519, 1521, 1528, 1535, 1536, 1630, 1632, 1727: oled_data = 16'b1111111000111011;
         2113, 2208, 2302, 2303, 2304, 2305, 2398, 2400, 2495, 3070: oled_data = 16'b1111111000111011;
         3072, 3167, 3168, 3169, 3263, 3648, 3743, 3744, 3838, 3840: oled_data = 16'b1111111000111011;
         3841, 3934, 3935, 3936, 4031, 4417, 4512, 4513, 4607, 4608: oled_data = 16'b1111111000111011;
         4702, 4703, 4704, 4705, 4798, 5184, 5279, 5280, 5281, 5375: oled_data = 16'b1111111000111011;
         5376, 5471, 5472, 5473, 5567, 6047, 6048, 6142: oled_data = 16'b1111111000111011;
         2, 4, 5, 10, 11, 18, 19, 26, 27, 29: oled_data = 16'b1111111011111101;
         34, 37, 42, 44, 45, 50, 51, 53, 58, 59: oled_data = 16'b1111111011111101;
         66, 67, 69, 74, 75, 77, 82, 83, 85, 90: oled_data = 16'b1111111011111101;
         92, 98, 106, 122, 138, 149, 154, 165, 173, 186: oled_data = 16'b1111111011111101;
         192, 199, 200, 201, 207, 208, 209, 214, 215, 223: oled_data = 16'b1111111011111101;
         224, 231, 233, 239, 240, 247, 248, 249, 255, 263: oled_data = 16'b1111111011111101;
         264, 271, 272, 279, 280, 281, 288, 303, 312, 329: oled_data = 16'b1111111011111101;
         344, 352, 353, 359, 361, 369, 383, 385, 391, 399: oled_data = 16'b1111111011111101;
         401, 407, 409, 415, 417, 423, 424, 431, 433, 439: oled_data = 16'b1111111011111101;
         440, 447, 449, 455, 465, 471, 472, 479, 480, 487: oled_data = 16'b1111111011111101;
         488, 495, 503, 504, 512, 519, 527, 528, 535, 537: oled_data = 16'b1111111011111101;
         543, 545, 551, 552, 559, 567, 569, 575, 579, 586: oled_data = 16'b1111111011111101;
         587, 589, 596, 612, 613, 618, 619, 621, 627, 634: oled_data = 16'b1111111011111101;
         635, 637, 643, 644, 645, 660, 666, 668, 674, 675: oled_data = 16'b1111111011111101;
         676, 684, 690, 691, 693, 698, 699, 701, 706, 707: oled_data = 16'b1111111011111101;
         716, 724, 732, 733, 738, 749, 754, 755, 763, 773: oled_data = 16'b1111111011111101;
         779, 781, 787, 789, 797, 804, 805, 810, 813, 819: oled_data = 16'b1111111011111101;
         821, 827, 834, 835, 836, 837, 842, 850, 852, 853: oled_data = 16'b1111111011111101;
         858, 860, 861, 866, 868, 874, 882, 890, 906, 914: oled_data = 16'b1111111011111101;
         917, 941, 947, 954, 960, 967, 968, 975, 976, 977: oled_data = 16'b1111111011111101;
         982, 984, 991, 992, 999, 1000, 1001, 1007, 1009, 1015: oled_data = 16'b1111111011111101;
         1016, 1023, 1024, 1025, 1040, 1047, 1048, 1049, 1056, 1064: oled_data = 16'b1111111011111101;
         1072, 1088, 1095, 1103, 1104, 1111, 1113, 1120, 1129, 1135: oled_data = 16'b1111111011111101;
         1137, 1144, 1151, 1159, 1161, 1167, 1169, 1176, 1183, 1185: oled_data = 16'b1111111011111101;
         1191, 1193, 1200, 1215, 1217, 1223, 1225, 1232, 1239, 1247: oled_data = 16'b1111111011111101;
         1248, 1255, 1256, 1263, 1265, 1271, 1272, 1279, 1280, 1287: oled_data = 16'b1111111011111101;
         1288, 1295, 1297, 1303, 1305, 1311, 1313, 1319, 1327, 1328: oled_data = 16'b1111111011111101;
         1336, 1343, 1346, 1347, 1354, 1355, 1362, 1370, 1372, 1378: oled_data = 16'b1111111011111101;
         1380, 1387, 1396, 1397, 1402, 1405, 1411, 1418, 1421, 1426: oled_data = 16'b1111111011111101;
         1435, 1437, 1442, 1444, 1445, 1450, 1453, 1458, 1461, 1475: oled_data = 16'b1111111011111101;
         1477, 1482, 1485, 1490, 1492, 1499, 1500, 1506, 1507, 1509: oled_data = 16'b1111111011111101;
         1515, 1517, 1523, 1525, 1530, 1531, 1533, 1539, 1628, 1634: oled_data = 16'b1111111011111101;
         1728, 1823, 1919, 1920, 2016, 2111, 2114, 2116, 2205, 2211: oled_data = 16'b1111111011111101;
         2307, 2308, 2396, 2402, 2496, 2591, 2593, 2687, 2688, 2784: oled_data = 16'b1111111011111101;
         2879, 2972, 2978, 2979, 3068, 3076, 3165, 3170, 3261, 3264: oled_data = 16'b1111111011111101;
         3359, 3361, 3456, 3551, 3552, 3647, 3650, 3740, 3746, 3747: oled_data = 16'b1111111011111101;
         3842, 3844, 3932, 3938, 3940, 4127, 4128, 4223, 4320, 4321: oled_data = 16'b1111111011111101;
         4414, 4415, 4514, 4516, 4604, 4605, 4610, 4612, 4701, 4796: oled_data = 16'b1111111011111101;
         4800, 4895, 4991, 4992, 5088, 5089, 5182, 5183, 5186, 5282: oled_data = 16'b1111111011111101;
         5283, 5284, 5372, 5373, 5378, 5380, 5469, 5476, 5568, 5663: oled_data = 16'b1111111011111101;
         5759, 5760, 5856, 5950, 5951, 5954, 6050, 6051, 6140: oled_data = 16'b1111111011111101;
         3, 12, 20, 28, 35, 43, 52, 61, 68, 76: oled_data = 16'b1111111100111101;
         84, 91, 99, 100, 101, 108, 109, 115, 116, 117: oled_data = 16'b1111111100111101;
         123, 124, 125, 131, 132, 133, 139, 141, 147, 148: oled_data = 16'b1111111100111101;
         156, 157, 162, 163, 170, 171, 172, 178, 180, 187: oled_data = 16'b1111111100111101;
         188, 189, 206, 222, 230, 238, 246, 254, 257, 262: oled_data = 16'b1111111100111101;
         270, 278, 286, 289, 294, 295, 296, 304, 305, 311: oled_data = 16'b1111111100111101;
         318, 327, 328, 334, 335, 337, 343, 351, 375, 376: oled_data = 16'b1111111100111101;
         377, 382, 384, 390, 393, 398, 400, 406, 408, 422: oled_data = 16'b1111111100111101;
         425, 432, 438, 441, 446, 448, 454, 456, 462, 464: oled_data = 16'b1111111100111101;
         470, 473, 478, 489, 494, 497, 518, 520, 526, 529: oled_data = 16'b1111111100111101;
         544, 553, 561, 566, 580, 588, 595, 597, 611, 659: oled_data = 16'b1111111100111101;
         661, 669, 683, 708, 715, 717, 725, 731, 739, 740: oled_data = 16'b1111111100111101;
         756, 764, 772, 780, 788, 796, 803, 811, 820, 828: oled_data = 16'b1111111100111101;
         844, 851, 859, 867, 869, 875, 877, 883, 884, 885: oled_data = 16'b1111111100111101;
         891, 892, 899, 900, 908, 909, 915, 916, 923, 924: oled_data = 16'b1111111100111101;
         925, 931, 932, 939, 940, 946, 948, 955, 957, 1006: oled_data = 16'b1111111100111101;
         1022, 1031, 1038, 1054, 1057, 1062, 1063, 1065, 1070, 1071: oled_data = 16'b1111111100111101;
         1073, 1078, 1081, 1086, 1087, 1089, 1094, 1096, 1105, 1110: oled_data = 16'b1111111100111101;
         1112, 1119, 1136, 1142, 1143, 1145, 1152, 1160, 1166, 1168: oled_data = 16'b1111111100111101;
         1174, 1175, 1177, 1184, 1192, 1199, 1207, 1209, 1214, 1216: oled_data = 16'b1111111100111101;
         1222, 1224, 1230, 1231, 1233, 1238, 1240, 1246, 1249, 1254: oled_data = 16'b1111111100111101;
         1264, 1270, 1278, 1286, 1289, 1294, 1296, 1304, 1312, 1318: oled_data = 16'b1111111100111101;
         1320, 1334, 1337, 1348, 1356, 1357, 1363, 1365, 1371, 1373: oled_data = 16'b1111111100111101;
         1379, 1389, 1395, 1403, 1404, 1413, 1419, 1427, 1428, 1436: oled_data = 16'b1111111100111101;
         1451, 1460, 1467, 1469, 1476, 1484, 1491, 1508, 1516, 1524: oled_data = 16'b1111111100111101;
         1540, 1629, 1635, 1724, 1729, 1824, 1918, 1921, 2014, 2015: oled_data = 16'b1111111100111101;
         2017, 2115, 2204, 2300, 2397, 2403, 2404, 2492, 2497, 2590: oled_data = 16'b1111111100111101;
         2592, 2782, 2783, 2785, 2883, 2973, 2980, 3075, 3164, 3172: oled_data = 16'b1111111100111101;
         3260, 3358, 3360, 3455, 3457, 3550, 3651, 3652, 3741, 3748: oled_data = 16'b1111111100111101;
         3836, 3939, 4028, 4033, 4222, 4224, 4225, 4319, 4419, 4420: oled_data = 16'b1111111100111101;
         4508, 4515, 4700, 4707, 4708, 4894, 4897, 4993, 5087, 5187: oled_data = 16'b1111111100111101;
         5188, 5277, 5379, 5468, 5475, 5564, 5569, 5662, 5664, 5761: oled_data = 16'b1111111100111101;
         5854, 5855, 5955, 5956, 6044, 6045, 6052: oled_data = 16'b1111111100111101;
         6, 30, 46, 54, 70, 78, 105, 110, 118, 129: oled_data = 16'b1111011001111011;
         134, 153, 158, 174, 590, 606, 622, 654, 694, 702: oled_data = 16'b1111011001111011;
         734, 750, 774, 822, 862, 865, 886, 889, 910, 913: oled_data = 16'b1111011001111011;
         918, 937, 942, 1350, 1398, 1406, 1414, 1478, 1518, 1534: oled_data = 16'b1111011001111011;
         1633, 2206, 2880, 2974, 2975, 2977, 3166, 4416, 4606, 5185: oled_data = 16'b1111011001111011;
         5470, 6046: oled_data = 16'b1111011001111011;
         13, 21, 36, 60, 93, 114, 130, 146, 193, 217: oled_data = 16'b1111011011111101;
         225, 232, 241, 256, 273, 287, 297, 319, 321, 367: oled_data = 16'b1111011011111101;
         392, 463, 486, 496, 502, 510, 521, 560, 578, 581: oled_data = 16'b1111011011111101;
         594, 603, 605, 610, 626, 628, 642, 650, 653, 658: oled_data = 16'b1111011011111101;
         682, 730, 741, 747, 757, 765, 786, 795, 812, 818: oled_data = 16'b1111011011111101;
         829, 845, 898, 938, 961, 974, 983, 985, 993, 1008: oled_data = 16'b1111011011111101;
         1017, 1030, 1032, 1033, 1039, 1055, 1127, 1153, 1208, 1321: oled_data = 16'b1111011011111101;
         1335, 1349, 1364, 1388, 1394, 1410, 1412, 1420, 1429, 1452: oled_data = 16'b1111011011111101;
         1459, 1468, 1483, 1498, 1522, 1825, 2301, 2306, 2493, 2882: oled_data = 16'b1111011011111101;
         2884, 3553, 3837, 4029, 4032, 4129, 4418, 4611, 4896, 5474: oled_data = 16'b1111011011111101;
         5565, 5665, 5857, 6141: oled_data = 16'b1111011011111101;
         25, 41, 65, 89, 96, 103, 112, 120, 127, 142: oled_data = 16'b1111011000111011;
         144, 151, 167, 169, 176, 177, 183, 190, 582, 584: oled_data = 16'b1111011000111011;
         599, 614, 624, 633, 640, 648, 662, 673, 679, 688: oled_data = 16'b1111011000111011;
         697, 704, 712, 718, 726, 728, 737, 745, 753, 760: oled_data = 16'b1111011000111011;
         767, 776, 793, 798, 801, 807, 816, 839, 841, 847: oled_data = 16'b1111011000111011;
         857, 870, 873, 880, 887, 895, 905, 920, 928, 935: oled_data = 16'b1111011000111011;
         945, 951, 1345, 1359, 1361, 1366, 1369, 1374, 1376, 1383: oled_data = 16'b1111011000111011;
         1385, 1392, 1401, 1408, 1417, 1433, 1447, 1449, 1455, 1463: oled_data = 16'b1111011000111011;
         1470, 1480, 1486, 1489, 1503, 1512, 1520, 1526, 1527, 1529: oled_data = 16'b1111011000111011;
         1537, 1631, 2112, 2207, 2209, 2399, 2401, 2881, 2976, 3071: oled_data = 16'b1111011000111011;
         3073, 3745, 3839, 3937, 4511, 4609, 4799, 5374, 5377, 5952: oled_data = 16'b1111011000111011;
         6049, 6143: oled_data = 16'b1111011000111011;
         94, 97, 113, 121, 126, 137, 145, 150, 166, 182: oled_data = 16'b1111111001111011;
         185, 630, 638, 646, 678, 742, 758, 766, 806, 814: oled_data = 16'b1111111001111011;
         838, 879, 881, 888, 894, 897, 904, 950, 953, 1390: oled_data = 16'b1111111001111011;
         1422, 1430, 1438, 1510, 2494, 3649, 3742, 4030, 4510, 5566: oled_data = 16'b1111111001111011;
         5953: oled_data = 16'b1111111001111011;
         107, 140, 155, 164, 179, 181, 198, 302, 310, 313: oled_data = 16'b1111011100111101;
         326, 342, 345, 350, 358, 360, 366, 374, 414, 416: oled_data = 16'b1111011100111101;
         430, 481, 505, 513, 534, 536, 542, 550, 558, 568: oled_data = 16'b1111011100111101;
         574, 604, 620, 636, 652, 667, 685, 692, 709, 723: oled_data = 16'b1111011100111101;
         771, 876, 893, 901, 907, 922, 930, 933, 949, 956: oled_data = 16'b1111011100111101;
         966, 969, 990, 998, 1014, 1046, 1080, 1097, 1102, 1118: oled_data = 16'b1111011100111101;
         1121, 1126, 1134, 1150, 1158, 1182, 1190, 1201, 1206, 1241: oled_data = 16'b1111011100111101;
         1257, 1262, 1281, 1302, 1310, 1326, 1329, 1342, 1381, 1443: oled_data = 16'b1111011100111101;
         1493, 1501, 1532, 1636, 1725, 1822, 2110, 2212, 2686, 2689: oled_data = 16'b1111011100111101;
         2878, 3069, 3171, 3265, 3454, 3646, 3843, 3933, 4126, 4318: oled_data = 16'b1111011100111101;
         4509, 4797, 4801, 4990, 5086, 5276, 5758: oled_data = 16'b1111011100111101;
         194, 202, 204, 210, 218, 242, 252, 261, 267, 276: oled_data = 16'b1111111110111110;
         285, 314, 346, 402, 410, 474, 482, 508, 514, 546: oled_data = 16'b1111111110111110;
         554, 557, 962, 970, 994, 1002, 1010, 1018, 1029, 1034: oled_data = 16'b1111111110111110;
         1042, 1082, 1210, 1234, 1242, 1258, 1266, 1285, 1298, 1308: oled_data = 16'b1111111110111110;
         1330, 1821, 1826, 2498, 2690, 2692, 2787, 3266, 3357, 3554: oled_data = 16'b1111111110111110;
         3556, 3645, 4034, 4130, 4322, 4412, 4898, 5092, 5180, 5570: oled_data = 16'b1111111110111110;
         5762, 5858: oled_data = 16'b1111111110111110;
         195, 197, 203, 205, 211, 213, 220, 228, 229, 236: oled_data = 16'b1111111110111111;
         237, 244, 253, 259, 269, 275, 277, 283, 338, 341: oled_data = 16'b1111111110111111;
         378, 386, 394, 418, 442, 453, 466, 498, 506, 522: oled_data = 16'b1111111110111111;
         525, 530, 533, 541, 573, 963, 965, 971, 972, 979: oled_data = 16'b1111111110111111;
         980, 987, 989, 995, 997, 1004, 1005, 1011, 1013, 1019: oled_data = 16'b1111111110111111;
         1020, 1021, 1026, 1027, 1036, 1044, 1045, 1051, 1052, 1053: oled_data = 16'b1111111110111111;
         1058, 1074, 1098, 1146, 1165, 1178, 1202, 1205, 1221, 1229: oled_data = 16'b1111111110111111;
         1250, 1261, 1274, 1282, 1290, 1309, 1322, 1332, 1333, 1338: oled_data = 16'b1111111110111111;
         1341, 1730, 1732, 1820, 1922, 2109, 2588, 2594, 2877, 3268: oled_data = 16'b1111111110111111;
         3362, 4125, 4802, 4994, 5085, 5661, 5859, 5948: oled_data = 16'b1111111110111111;
         196, 245, 381, 411, 450, 500, 532, 981, 1069, 1114: oled_data = 16'b1111011111111111;
         1212, 1235, 1237, 2691: oled_data = 16'b1111011111111111;
         212, 219, 235, 243, 251, 260, 268, 284, 291, 292: oled_data = 16'b1111111111111111;
         293, 299, 300, 301, 307, 308, 309, 315, 316, 317: oled_data = 16'b1111111111111111;
         323, 324, 325, 330, 331, 332, 333, 339, 340, 347: oled_data = 16'b1111111111111111;
         348, 349, 355, 356, 357, 363, 364, 365, 371, 372: oled_data = 16'b1111111111111111;
         373, 379, 380, 387, 388, 395, 396, 397, 403, 404: oled_data = 16'b1111111111111111;
         405, 412, 413, 419, 420, 421, 427, 428, 435, 436: oled_data = 16'b1111111111111111;
         443, 444, 445, 451, 452, 459, 460, 467, 468, 469: oled_data = 16'b1111111111111111;
         475, 476, 477, 483, 485, 491, 492, 499, 507, 515: oled_data = 16'b1111111111111111;
         516, 523, 524, 539, 540, 547, 548, 549, 555, 563: oled_data = 16'b1111111111111111;
         564, 571, 572, 964, 973, 988, 996, 1003, 1012, 1028: oled_data = 16'b1111111111111111;
         1035, 1037, 1043, 1059, 1060, 1061, 1067, 1068, 1075, 1076: oled_data = 16'b1111111111111111;
         1077, 1083, 1084, 1085, 1091, 1092, 1093, 1099, 1100, 1101: oled_data = 16'b1111111111111111;
         1106, 1107, 1108, 1109, 1115, 1116, 1123, 1124, 1125, 1130: oled_data = 16'b1111111111111111;
         1131, 1132, 1133, 1139, 1140, 1141, 1147, 1148, 1149, 1155: oled_data = 16'b1111111111111111;
         1156, 1157, 1162, 1163, 1171, 1172, 1173, 1179, 1180, 1181: oled_data = 16'b1111111111111111;
         1187, 1189, 1195, 1196, 1197, 1203, 1204, 1211, 1213, 1219: oled_data = 16'b1111111111111111;
         1220, 1227, 1228, 1243, 1244, 1251, 1252, 1253, 1259, 1260: oled_data = 16'b1111111111111111;
         1267, 1268, 1275, 1276, 1277, 1283, 1284, 1291, 1292, 1299: oled_data = 16'b1111111111111111;
         1300, 1306, 1307, 1315, 1316, 1323, 1324, 1325, 1331, 1339: oled_data = 16'b1111111111111111;
         1731, 1827, 1828, 1916, 1917, 1923, 1924, 2013, 2019, 2020: oled_data = 16'b1111111111111111;
         2108, 2499, 2589, 2595, 2684, 2685, 2780, 2781, 2788, 3267: oled_data = 16'b1111111111111111;
         3356, 3363, 3364, 3452, 3453, 3458, 3459, 3460, 3548, 3549: oled_data = 16'b1111111111111111;
         3555, 3644, 4035, 4036, 4124, 4131, 4132, 4220, 4221, 4227: oled_data = 16'b1111111111111111;
         4228, 4316, 4317, 4413, 4803, 4804, 4892, 4893, 4899, 4900: oled_data = 16'b1111111111111111;
         4988, 4989, 4995, 4996, 5084, 5091, 5571, 5572, 5660, 5666: oled_data = 16'b1111111111111111;
         5667, 5668, 5756, 5757, 5763, 5764, 5852, 5853, 5860: oled_data = 16'b1111111111111111;
         216, 265, 457, 602, 677, 722, 746, 770, 778, 802: oled_data = 16'b1111111011111100;
         826, 1386, 1434, 1466, 1514, 1538, 2210, 3074: oled_data = 16'b1111111011111100;
         221, 258, 266, 306, 458, 493, 556, 565, 570, 1090: oled_data = 16'b1111011110111111;
         1138, 1218, 4226, 4324: oled_data = 16'b1111011110111111;
         226: oled_data = 16'b1111111101111110;
         227, 234, 250, 274, 282, 290, 426, 434, 461, 484: oled_data = 16'b1111011110111110;
         490, 562, 978, 986, 1050, 1066, 1188, 1269, 1293, 1317: oled_data = 16'b1111011110111110;
         2018, 2500, 2596, 2786, 5090, 5949: oled_data = 16'b1111011110111110;
         298, 322, 354, 362, 370, 389, 429, 437, 501, 509: oled_data = 16'b1111111111111110;
         531, 538, 1117, 1122, 1154, 1186, 1226, 1236, 1245, 1301: oled_data = 16'b1111111111111110;
         1314, 2876, 4323: oled_data = 16'b1111111111111110;
         320, 368, 700, 1273: oled_data = 16'b1111011100111100;
         336, 511, 629, 651, 714, 762, 794, 843, 1041, 1079: oled_data = 16'b1111011011111100;
         1198, 1474, 1541, 4706: oled_data = 16'b1111011011111100;
         517, 1164, 1170, 1194, 1340, 2012, 5181: oled_data = 16'b1111011111111110;
         748, 1128: oled_data = 16'b1111111100111100;
         878: oled_data = 16'b1111011000111100;
         902: oled_data = 16'b1111111000111100;
         926, 3262: oled_data = 16'b1111011001111100;
         934, 1726, 5278: oled_data = 16'b1111111001111100;
         1542: oled_data = 16'b0011100110000110;
         1543, 1545, 1547, 1549, 1551, 1553, 1556, 1558, 1559, 1561: oled_data = 16'b0001000010000010;
         1562, 1564, 1566, 1568, 1569, 1570, 1572, 1573, 1574, 1576: oled_data = 16'b0001000010000010;
         1578, 1581, 1582, 1584, 1586, 1588, 1590, 1591, 1592, 1595: oled_data = 16'b0001000010000010;
         1597, 1599, 1601, 1603, 1605, 1606, 1609, 1610, 1612, 1616: oled_data = 16'b0001000010000010;
         1618, 1620, 1622, 1623, 1625, 1638, 1640, 1641, 1643, 1645: oled_data = 16'b0001000010000010;
         1646, 1650, 1653, 1655, 1656, 1660, 1662, 1663, 1666, 1673: oled_data = 16'b0001000010000010;
         1675, 1678, 1679, 1682, 1685, 1689, 1690, 1692, 1694, 1695: oled_data = 16'b0001000010000010;
         1697, 1698, 1702, 1704, 1706, 1708, 1710, 1711, 1714, 1717: oled_data = 16'b0001000010000010;
         1719, 1721, 1734, 1735, 1736, 1817, 1818, 1831, 1926, 2009: oled_data = 16'b0001000010000010;
         2023, 2106, 2118, 2129, 2130, 2191, 2193, 2201, 2215, 2222: oled_data = 16'b0001000010000010;
         2225, 2226, 2285, 2286, 2288, 2289, 2290, 2298, 2310, 2319: oled_data = 16'b0001000010000010;
         2322, 2323, 2382, 2387, 2393, 2407, 2477, 2478, 2483, 2489: oled_data = 16'b0001000010000010;
         2502, 2509, 2510, 2515, 2572, 2574, 2578, 2586, 2598, 2606: oled_data = 16'b0001000010000010;
         2607, 2610, 2612, 2669, 2670, 2673, 2675, 2681, 2695, 2703: oled_data = 16'b0001000010000010;
         2704, 2706, 2765, 2767, 2769, 2770, 2778, 2790, 2799, 2801: oled_data = 16'b0001000010000010;
         2802, 2864, 2873, 2887, 3065, 3079, 3162, 3174, 3257, 3270: oled_data = 16'b0001000010000010;
         3271, 3272, 3273, 3274, 3275, 3276, 3277, 3278, 3279, 3280: oled_data = 16'b0001000010000010;
         3281, 3282, 3283, 3285, 3286, 3287, 3288, 3289, 3290, 3291: oled_data = 16'b0001000010000010;
         3292, 3293, 3294, 3295, 3297, 3298, 3299, 3301, 3303, 3304: oled_data = 16'b0001000010000010;
         3305, 3306, 3307, 3308, 3309, 3310, 3312, 3314, 3316, 3317: oled_data = 16'b0001000010000010;
         3318, 3319, 3320, 3321, 3322, 3323, 3324, 3325, 3326, 3327: oled_data = 16'b0001000010000010;
         3328, 3329, 3330, 3331, 3333, 3335, 3336, 3337, 3339, 3341: oled_data = 16'b0001000010000010;
         3342, 3343, 3344, 3346, 3348, 3349, 3350, 3352, 3354, 3366: oled_data = 16'b0001000010000010;
         3369, 3372, 3375, 3378, 3380, 3383, 3386, 3388, 3391, 3393: oled_data = 16'b0001000010000010;
         3395, 3397, 3398, 3400, 3403, 3406, 3407, 3409, 3410, 3412: oled_data = 16'b0001000010000010;
         3415, 3418, 3420, 3423, 3426, 3428, 3430, 3432, 3434, 3436: oled_data = 16'b0001000010000010;
         3438, 3440, 3442, 3443, 3445, 3447, 3449, 3450, 3463, 3559: oled_data = 16'b0001000010000010;
         3641, 3654, 3737, 3750, 3758, 3760, 3762, 3764, 3765, 3768: oled_data = 16'b0001000010000010;
         3770, 3772, 3776, 3778, 3779, 3781, 3782, 3784, 3787, 3788: oled_data = 16'b0001000010000010;
         3790, 3792, 3794, 3796, 3798, 3800, 3801, 3802, 3805, 3806: oled_data = 16'b0001000010000010;
         3808, 3809, 3811, 3813, 3815, 3818, 3820, 3821, 3822, 3824: oled_data = 16'b0001000010000010;
         3825, 3827, 3834, 3847, 3854, 3856, 3857, 3859, 3863, 3865: oled_data = 16'b0001000010000010;
         3867, 3870, 3871, 3875, 3877, 3879, 3881, 3888, 3890, 3893: oled_data = 16'b0001000010000010;
         3894, 3899, 3900, 3902, 3903, 3905, 3908, 3910, 3913, 3915: oled_data = 16'b0001000010000010;
         3919, 3921, 3923, 3930, 3942, 4025, 4038, 4121, 4122, 4218: oled_data = 16'b0001000010000010;
         4230, 4313, 4326, 4327, 4409, 4410, 4423, 4505, 4518, 4602: oled_data = 16'b0001000010000010;
         4615, 4697, 4698, 4710, 4806, 4889, 4890, 4903, 4914, 4915: oled_data = 16'b0001000010000010;
         4916, 4917, 4918, 4919, 4921, 4922, 4924, 4925, 4927, 4928: oled_data = 16'b0001000010000010;
         4929, 4930, 4931, 4933, 4935, 4936, 4937, 4939, 4940, 4941: oled_data = 16'b0001000010000010;
         4942, 4944, 4946, 4947, 4949, 4951, 4952, 4954, 4955, 4957: oled_data = 16'b0001000010000010;
         4959, 4960, 4962, 4963, 4964, 4965, 4966, 4967, 4968, 4969: oled_data = 16'b0001000010000010;
         4971, 4972, 4974, 4986, 4999, 5013, 5015, 5017, 5019, 5021: oled_data = 16'b0001000010000010;
         5027, 5028, 5030, 5033, 5034, 5036, 5039, 5041, 5043, 5046: oled_data = 16'b0001000010000010;
         5050, 5052, 5054, 5057, 5060, 5063, 5066, 5070, 5081, 5095: oled_data = 16'b0001000010000010;
         5106, 5166, 5178, 5190, 5202, 5203, 5263, 5273, 5286, 5358: oled_data = 16'b0001000010000010;
         5369, 5370, 5383, 5394, 5395, 5466, 5478, 5491, 5551, 5561: oled_data = 16'b0001000010000010;
         5574, 5575, 5646, 5657, 5658, 5671, 5682, 5742, 5753, 5767: oled_data = 16'b0001000010000010;
         5778, 5779, 5839, 5849, 5862, 5875, 5934, 5945, 5958, 5959: oled_data = 16'b0001000010000010;
         5970, 6031, 6042, 6055, 6067, 6127, 6138: oled_data = 16'b0001000010000010;
         1544, 1546, 1548, 1550, 1552, 1554, 1555, 1557, 1560, 1563: oled_data = 16'b0001000010000001;
         1565, 1567, 1571, 1575, 1577, 1579, 1580, 1583, 1585, 1587: oled_data = 16'b0001000010000001;
         1589, 1593, 1594, 1596, 1598, 1600, 1602, 1604, 1608, 1611: oled_data = 16'b0001000010000001;
         1613, 1615, 1617, 1619, 1621, 1624, 1639, 1644, 1647, 1649: oled_data = 16'b0001000010000001;
         1652, 1654, 1657, 1659, 1664, 1665, 1667, 1669, 1671, 1674: oled_data = 16'b0001000010000001;
         1677, 1680, 1683, 1686, 1688, 1691, 1699, 1701, 1703, 1705: oled_data = 16'b0001000010000001;
         1709, 1712, 1715, 1718, 1722, 1830, 1913, 2010, 2022, 2105: oled_data = 16'b0001000010000001;
         2119, 2128, 2192, 2202, 2223, 2227, 2287, 2297, 2311, 2318: oled_data = 16'b0001000010000001;
         2324, 2381, 2386, 2394, 2406, 2413, 2419, 2476, 2482, 2503: oled_data = 16'b0001000010000001;
         2516, 2585, 2611, 2674, 2682, 2694, 2705, 2707, 2766, 2768: oled_data = 16'b0001000010000001;
         2777, 2791, 2800, 2863, 2874, 2886, 2969, 2983, 3066, 3078: oled_data = 16'b0001000010000001;
         3161, 3175, 3258, 3284, 3296, 3300, 3302, 3311, 3313, 3315: oled_data = 16'b0001000010000001;
         3332, 3334, 3338, 3340, 3345, 3347, 3351, 3368, 3370, 3371: oled_data = 16'b0001000010000001;
         3373, 3374, 3376, 3377, 3379, 3381, 3382, 3384, 3385, 3387: oled_data = 16'b0001000010000001;
         3389, 3390, 3392, 3394, 3396, 3399, 3401, 3402, 3404, 3408: oled_data = 16'b0001000010000001;
         3411, 3413, 3414, 3416, 3417, 3419, 3421, 3422, 3424, 3425: oled_data = 16'b0001000010000001;
         3427, 3429, 3431, 3433, 3435, 3439, 3441, 3444, 3446, 3448: oled_data = 16'b0001000010000001;
         3462, 3545, 3558, 3642, 3655, 3738, 3751, 3759, 3761, 3766: oled_data = 16'b0001000010000001;
         3769, 3771, 3773, 3775, 3777, 3783, 3786, 3789, 3791, 3795: oled_data = 16'b0001000010000001;
         3799, 3804, 3810, 3814, 3816, 3819, 3823, 3826, 3846, 3853: oled_data = 16'b0001000010000001;
         3858, 3860, 3862, 3864, 3869, 3872, 3874, 3876, 3880, 3882: oled_data = 16'b0001000010000001;
         3884, 3886, 3889, 3892, 3895, 3897, 3898, 3904, 3907, 3909: oled_data = 16'b0001000010000001;
         3912, 3914, 3917, 3922, 3929, 3943, 4026, 4039, 4134, 4231: oled_data = 16'b0001000010000001;
         4314, 4422, 4519, 4601, 4711, 4794, 4807, 4902, 4920, 4923: oled_data = 16'b0001000010000001;
         4932, 4938, 4945, 4948, 4950, 4953, 4956, 4958, 4961, 4970: oled_data = 16'b0001000010000001;
         4973, 4975, 4985, 4998, 5010, 5012, 5020, 5022, 5023, 5025: oled_data = 16'b0001000010000001;
         5029, 5031, 5038, 5040, 5044, 5047, 5049, 5055, 5058, 5061: oled_data = 16'b0001000010000001;
         5064, 5067, 5069, 5107, 5167, 5177, 5191, 5262, 5274, 5287: oled_data = 16'b0001000010000001;
         5298, 5299, 5359, 5382, 5455, 5490, 5550, 5562, 5587, 5647: oled_data = 16'b0001000010000001;
         5670, 5683, 5743, 5766, 5850, 5863, 5874, 5935, 5946, 6030: oled_data = 16'b0001000010000001;
         6054, 6066, 6126, 6137: oled_data = 16'b0001000010000001;
         1607, 1614, 1648, 1651, 1658, 1668, 1670, 1672, 1676, 1681: oled_data = 16'b0001000001000010;
         1684, 1687, 1700, 1713, 1716, 1914, 2224, 2385, 2414, 2420: oled_data = 16'b0001000001000010;
         2490, 2599, 2970, 2982, 3546, 3767, 3774, 3785, 3803, 3817: oled_data = 16'b0001000001000010;
         3833, 3861, 3868, 3873, 3883, 3885, 3887, 3891, 3896, 3906: oled_data = 16'b0001000001000010;
         3911, 3918, 4135, 4793, 4926, 4934, 4943, 5011, 5024, 5045: oled_data = 16'b0001000001000010;
         5048, 5056, 5065, 5068, 5071, 5454, 5586, 6041: oled_data = 16'b0001000001000010;
         1626, 1742, 1756, 1758, 1772, 1774, 1781, 1793, 1802, 1806: oled_data = 16'b0010000011000011;
         1809, 2321: oled_data = 16'b0010000011000011;
         1627: oled_data = 16'b1011010100110101;
         1637, 2117, 2213, 2981, 3173, 3845, 4613, 5189, 5477: oled_data = 16'b1101010111111000;
         1642, 1661, 1693, 1696, 1707, 1720, 1927, 2214, 2573, 2579: oled_data = 16'b0001000001000001;
         2702, 2865, 3353, 3367, 3405, 3437, 3763, 3780, 3793, 3797: oled_data = 16'b0001000001000001;
         3807, 3812, 3855, 3866, 3878, 3901, 3916, 3920, 4217, 4506: oled_data = 16'b0001000001000001;
         4614, 5014, 5016, 5018, 5026, 5032, 5035, 5037, 5042, 5051: oled_data = 16'b0001000001000001;
         5053, 5059, 5062, 5082, 5094, 5465, 5479, 5754, 5838, 5971: oled_data = 16'b0001000001000001;
         1723, 2395, 2491, 2971, 3067, 3739, 3931, 4507, 4603, 4795: oled_data = 16'b0111001101001101;
         5371, 5563, 6043: oled_data = 16'b0111001101001101;
         1733, 2501, 2789, 4037, 4229, 4325, 4805, 5861: oled_data = 16'b1101011001111001;
         1737, 1739, 1763, 1766, 1768, 1778, 1790, 1812: oled_data = 16'b0010000100000011;
         1738, 1740, 1762, 1767, 1779, 1791, 1794, 1796, 1801, 1811: oled_data = 16'b0001100011000100;
         4019: oled_data = 16'b0001100011000100;
         1741, 1744, 1746, 1749, 1751, 1752, 1754, 1761, 1764, 1769: oled_data = 16'b0001100011000011;
         1775, 1777, 1783, 1786, 1787, 1789, 1798, 1804, 1807, 1813: oled_data = 16'b0001100011000011;
         1816, 2608, 2671, 2862, 3176, 3757, 3950, 3952, 3953, 3954: oled_data = 16'b0001100011000011;
         3955, 3956, 3958, 3959, 3960, 3961, 3963, 3964, 3965, 3966: oled_data = 16'b0001100011000011;
         3967, 3968, 3969, 3970, 3971, 3972, 3973, 3975, 3976, 3977: oled_data = 16'b0001100011000011;
         3978, 3980, 3981, 3983, 3984, 3985, 3986, 3988, 3989, 3990: oled_data = 16'b0001100011000011;
         3991, 3992, 3993, 3994, 3995, 3996, 3998, 3999, 4000, 4001: oled_data = 16'b0001100011000011;
         4002, 4003, 4004, 4005, 4006, 4007, 4008, 4009, 4010, 4011: oled_data = 16'b0001100011000011;
         4012, 4014, 4015, 4017, 4018, 4913, 5009, 5297, 5489, 5681: oled_data = 16'b0001100011000011;
         5969, 6065: oled_data = 16'b0001100011000011;
         1743, 1755, 1757, 1765, 1773, 1782, 1803, 1805, 1808: oled_data = 16'b0001100100000100;
         1745, 1750, 1753, 1776, 1788, 2127, 2190, 2317, 2418, 2605: oled_data = 16'b0010000100000100;
         2609, 2672, 3464, 3560, 3848, 4328, 4424, 4616, 4818, 4819: oled_data = 16'b0010000100000100;
         4820, 4821, 4822, 4823, 4824, 4825, 4826, 4827, 4828, 4829: oled_data = 16'b0010000100000100;
         4830, 4831, 4832, 4833, 4834, 4835, 4836, 4837, 4838, 4839: oled_data = 16'b0010000100000100;
         4840, 4841, 4842, 4843, 4844, 4845, 4846, 4847, 4848, 4849: oled_data = 16'b0010000100000100;
         4850, 4851, 4852, 4853, 4854, 4855, 4856, 4857, 4858, 4859: oled_data = 16'b0010000100000100;
         4860, 4861, 4862, 4863, 4864, 4865, 4866, 4867, 4868, 4869: oled_data = 16'b0010000100000100;
         4870, 4871, 4872, 4873, 4874, 4875, 4876, 4877, 4878, 4904: oled_data = 16'b0010000100000100;
         5000, 5384, 5576, 5672, 5768, 5960, 6056: oled_data = 16'b0010000100000100;
         1747, 1759, 1771, 1780, 1784, 1792, 1795, 1797, 1800, 1810: oled_data = 16'b0001100100000011;
         1815, 2384, 3951, 3957, 3962, 3974, 3979, 3982, 3987, 3997: oled_data = 16'b0001100100000011;
         4013, 4016: oled_data = 16'b0001100100000011;
         1748, 1760, 1770, 1785, 1799, 1814: oled_data = 16'b0010000011000100;
         1819, 1915, 2011, 2107, 2587, 2683, 2779, 2875, 3355, 3451: oled_data = 16'b0111001110001110;
         3547, 3643, 4123, 4219, 4315, 4411, 4891, 4987, 5083, 5179: oled_data = 16'b0111001110001110;
         5659, 5755, 5851, 5947: oled_data = 16'b0111001110001110;
         1829, 2693, 3461, 4133, 4901, 5093: oled_data = 16'b1100111010111010;
         1832, 2194, 3661, 4080, 4085, 4119, 4148, 4154, 4161, 4170: oled_data = 16'b0100001000001000;
         4174, 4179, 4194, 4200, 4237, 4273, 4331, 4335, 4344, 4351: oled_data = 16'b0100001000001000;
         4354, 4357, 4360, 4363, 4367, 4383, 4386, 4389, 4392, 4394: oled_data = 16'b0100001000001000;
         4407, 4445, 4461, 4467, 4470, 4473, 4501, 4528, 4531, 4534: oled_data = 16'b0100001000001000;
         4537, 4544, 4547, 4550, 4552, 4555, 4561, 4577, 4582, 4585: oled_data = 16'b0100001000001000;
         4655, 4660, 4663, 4715, 4727, 4743, 4749, 4761, 4767, 4785: oled_data = 16'b0100001000001000;
         4908, 4911, 5077, 5101, 5104, 5171, 5270, 5363, 5487, 5555: oled_data = 16'b0100001000001000;
         5558, 5674, 5677, 5747, 5750, 5775, 5866, 5869, 5939, 6058: oled_data = 16'b0100001000001000;
         1833, 1841, 1963, 1996, 2034, 2094, 2097, 2103, 2132, 2571: oled_data = 16'b0111001111010000;
         2604, 2614, 2698, 2804, 2867, 2895, 2958, 2993, 3097, 3103: oled_data = 16'b0111001111010000;
         3123, 3136, 3147, 5108, 5122, 5131, 5147: oled_data = 16'b0111001111010000;
         1834, 1837, 1840, 1842, 1844, 1847, 1854, 1859, 1864, 1868: oled_data = 16'b0111110000010001;
         1873, 1877, 1880, 1883, 1889, 1905, 1945, 1947, 1957, 1966: oled_data = 16'b0111110000010001;
         1971, 1980, 1987, 1991, 1993, 1995, 1997, 2003, 2025, 2036: oled_data = 16'b0111110000010001;
         2093, 2102, 2133, 2188, 2196, 2217, 2295, 2316, 2377, 2505: oled_data = 16'b0111110000010001;
         2518, 2568, 2570, 2602, 2603, 2678, 2700, 2709, 2763, 2772: oled_data = 16'b0111110000010001;
         2775, 2793, 2794, 2891, 2894, 2900, 2902, 2907, 2923, 2936: oled_data = 16'b0111110000010001;
         2946, 2952, 2955, 2985, 2989, 2994, 2999, 3001, 3008, 3010: oled_data = 16'b0111110000010001;
         3013, 3017, 3022, 3025, 3028, 3034, 3038, 3040, 3044, 3046: oled_data = 16'b0111110000010001;
         3051, 3053, 3055, 3058, 3082, 3088, 3098, 3102, 3105, 3110: oled_data = 16'b0111110000010001;
         3113, 3122, 3128, 3135, 3137, 3145, 3148, 3159, 5114, 5121: oled_data = 16'b0111110000010001;
         5127, 5130, 5132, 5140, 5146, 5148: oled_data = 16'b0111110000010001;
         1835, 1836, 1839, 1843, 1848, 1850, 1852, 1853, 1856, 1857: oled_data = 16'b0111110000010000;
         1858, 1860, 1862, 1863, 1865, 1866, 1867, 1870, 1871, 1872: oled_data = 16'b0111110000010000;
         1875, 1876, 1879, 1881, 1882, 1884, 1885, 1887, 1888, 1890: oled_data = 16'b0111110000010000;
         1891, 1892, 1894, 1895, 1897, 1899, 1900, 1903, 1904, 1907: oled_data = 16'b0111110000010000;
         1909, 1910, 1929, 1935, 1937, 1938, 1940, 1942, 1948, 1950: oled_data = 16'b0111110000010000;
         1951, 1953, 1955, 1958, 1960, 1962, 1964, 1965, 1970, 1973: oled_data = 16'b0111110000010000;
         1974, 1976, 1978, 1982, 1983, 1985, 1989, 1990, 1992, 1998: oled_data = 16'b0111110000010000;
         2006, 2007, 2026, 2029, 2030, 2035, 2039, 2089, 2092, 2098: oled_data = 16'b0111110000010000;
         2121, 2123, 2124, 2134, 2184, 2186, 2197, 2199, 2218, 2229: oled_data = 16'b0111110000010000;
         2231, 2280, 2281, 2283, 2292, 2294, 2315, 2327, 2378, 2389: oled_data = 16'b0111110000010000;
         2391, 2409, 2423, 2472, 2473, 2486, 2487, 2519, 2581, 2583: oled_data = 16'b0111110000010000;
         2615, 2664, 2665, 2666, 2697, 2699, 2710, 2760, 2805, 2807: oled_data = 16'b0111110000010000;
         2856, 2857, 2859, 2860, 2868, 2871, 2892, 2899, 2901, 2904: oled_data = 16'b0111110000010000;
         2906, 2909, 2910, 2912, 2913, 2915, 2916, 2918, 2919, 2921: oled_data = 16'b0111110000010000;
         2922, 2924, 2925, 2927, 2928, 2930, 2931, 2933, 2935, 2937: oled_data = 16'b0111110000010000;
         2939, 2940, 2942, 2943, 2944, 2947, 2949, 2950, 2957, 2962: oled_data = 16'b0111110000010000;
         2964, 2966, 2991, 2992, 2995, 2997, 3002, 3004, 3005, 3007: oled_data = 16'b0111110000010000;
         3011, 3014, 3016, 3019, 3021, 3024, 3027, 3029, 3030, 3032: oled_data = 16'b0111110000010000;
         3035, 3037, 3041, 3043, 3047, 3048, 3060, 3062, 3081, 3085: oled_data = 16'b0111110000010000;
         3089, 3091, 3092, 3094, 3096, 3099, 3101, 3104, 3108, 3116: oled_data = 16'b0111110000010000;
         3118, 3124, 3127, 3131, 3134, 3138, 3141, 3146, 3151, 3153: oled_data = 16'b0111110000010000;
         3156, 5110, 5112, 5119, 5137, 5143: oled_data = 16'b0111110000010000;
         1838, 1845, 1849, 1931, 1933, 2000, 2002, 2037, 2090, 2100: oled_data = 16'b0111010000010000;
         2187, 2195, 2220, 2326, 2411, 2475, 2506, 2679, 2762, 2773: oled_data = 16'b0111010000010000;
         2796, 2870, 2890, 2893, 2903, 3049, 3052, 3056, 3059, 3063: oled_data = 16'b0111010000010000;
         3111, 3114, 3121, 3129, 3132, 3140, 3143, 3154, 5154: oled_data = 16'b0111010000010000;
         1846, 1851, 1855, 1861, 1869, 1874, 1878, 1896, 1901, 1906: oled_data = 16'b0111101111010000;
         1944, 1946, 1956, 1959, 1967, 1969, 1972, 1977, 1979, 1981: oled_data = 16'b0111101111010000;
         1986, 1988, 1994, 2004, 2027, 2038, 2088, 2101, 2313, 2376: oled_data = 16'b0111101111010000;
         2474, 2507, 2569, 2601, 2667, 2677, 2774, 2795, 2858, 2889: oled_data = 16'b0111101111010000;
         2905, 2908, 2911, 2914, 2917, 2920, 2926, 2929, 2932, 2934: oled_data = 16'b0111101111010000;
         2938, 2941, 2945, 2948, 2951, 2953, 2956, 2986, 2988, 2990: oled_data = 16'b0111101111010000;
         2998, 3000, 3003, 3009, 3012, 3018, 3020, 3023, 3026, 3031: oled_data = 16'b0111101111010000;
         3033, 3039, 3042, 3045, 3050, 3054, 3057, 3083, 3087, 3106: oled_data = 16'b0111101111010000;
         3109, 3112, 3120, 3149, 3158, 5115, 5117, 5124, 5126, 5129: oled_data = 16'b0111101111010000;
         5133, 5135, 5139, 5141, 5145, 5150, 5152, 5156, 5159, 5161: oled_data = 16'b0111101111010000;
         5162, 5164: oled_data = 16'b0111101111010000;
         1886, 1893, 1911, 1930, 1932, 1934, 1936, 1941, 1949, 1952: oled_data = 16'b0111101111010001;
         1954, 1961, 1975, 1984, 1999, 2001, 2091, 2099, 2125, 2185: oled_data = 16'b0111101111010001;
         2219, 2230, 2282, 2293, 2410, 2422, 2711, 2761, 2797, 2869: oled_data = 16'b0111101111010001;
         2963, 2967, 3006, 3015, 3036, 3061, 3115, 3125, 3130, 3133: oled_data = 16'b0111101111010001;
         3139, 3142, 3144, 3152, 3155, 5109, 5111, 5113, 5116, 5118: oled_data = 16'b0111101111010001;
         5120, 5123, 5136, 5138, 5142, 5144, 5149, 5153, 5155, 5158: oled_data = 16'b0111101111010001;
         1898, 1902, 1908, 1943, 1968, 2005, 2028, 2314, 2485, 2954: oled_data = 16'b0111010000010001;
         2965, 2987, 3084, 3086, 3095, 3107, 3119, 3126, 3150, 3157: oled_data = 16'b0111010000010001;
         5134, 5151, 5157, 5160, 5163: oled_data = 16'b0111010000010001;
         1912, 2200: oled_data = 16'b0110001110001110;
         1925, 3365: oled_data = 16'b1101011010111001;
         1928, 2024, 2216, 2312, 2480, 2504, 2512, 2575, 2600, 2696: oled_data = 16'b0011101000001000;
         2888, 2984, 3563, 3566, 3569, 3573, 3575, 3580, 3582, 3584: oled_data = 16'b0011101000001000;
         3586, 3590, 3592, 3594, 3596, 3600, 3604, 3608, 3609, 3613: oled_data = 16'b0011101000001000;
         3615, 3619, 3621, 3623, 3625, 3627, 3629, 3631, 3636, 3639: oled_data = 16'b0011101000001000;
         3657, 3660, 3732, 3733, 3734, 3753, 3754, 3831, 3925, 3927: oled_data = 16'b0011101000001000;
         3945, 3946, 3947, 3948, 4022, 4041, 4045, 4048, 4050, 4054: oled_data = 16'b0011101000001000;
         4056, 4060, 4061, 4063, 4065, 4067, 4069, 4071, 4073, 4077: oled_data = 16'b0011101000001000;
         4079, 4082, 4086, 4088, 4090, 4092, 4095, 4096, 4098, 4100: oled_data = 16'b0011101000001000;
         4102, 4103, 4105, 4107, 4111, 4114, 4115, 4117, 4138, 4140: oled_data = 16'b0011101000001000;
         4143, 4147, 4150, 4152, 4155, 4157, 4159, 4163, 4165, 4166: oled_data = 16'b0011101000001000;
         4168, 4171, 4173, 4176, 4183, 4185, 4187, 4189, 4190, 4196: oled_data = 16'b0011101000001000;
         4202, 4204, 4205, 4208, 4210, 4212, 4214, 4233, 4234, 4238: oled_data = 16'b0011101000001000;
         4240, 4241, 4245, 4247, 4249, 4251, 4252, 4255, 4259, 4261: oled_data = 16'b0011101000001000;
         4263, 4269, 4271, 4275, 4276, 4277, 4280, 4282, 4283, 4284: oled_data = 16'b0011101000001000;
         4287, 4289, 4291, 4293, 4294, 4295, 4297, 4299, 4301, 4302: oled_data = 16'b0011101000001000;
         4304, 4307, 4308, 4310, 4311, 4329, 4337, 4339, 4340, 4342: oled_data = 16'b0011101000001000;
         4346, 4349, 4353, 4356, 4358, 4361, 4364, 4366, 4369, 4375: oled_data = 16'b0011101000001000;
         4377, 4381, 4388, 4391, 4396, 4398, 4401, 4405, 4426, 4428: oled_data = 16'b0011101000001000;
         4429, 4431, 4432, 4434, 4438, 4442, 4447, 4451, 4453, 4455: oled_data = 16'b0011101000001000;
         4457, 4464, 4466, 4469, 4475, 4478, 4480, 4484, 4486, 4488: oled_data = 16'b0011101000001000;
         4492, 4493, 4495, 4498, 4499, 4502, 4521, 4523, 4526, 4529: oled_data = 16'b0011101000001000;
         4532, 4536, 4539, 4540, 4542, 4545, 4548, 4551, 4554, 4557: oled_data = 16'b0011101000001000;
         4560, 4564, 4566, 4567, 4570, 4572, 4575, 4578, 4581, 4583: oled_data = 16'b0011101000001000;
         4586, 4591, 4593, 4599, 4618, 4620, 4622, 4623, 4626, 4628: oled_data = 16'b0011101000001000;
         4630, 4634, 4636, 4637, 4642, 4644, 4645, 4650, 4652, 4657: oled_data = 16'b0011101000001000;
         4658, 4661, 4664, 4666, 4668, 4670, 4672, 4674, 4675, 4680: oled_data = 16'b0011101000001000;
         4682, 4683, 4684, 4685, 4687, 4690, 4691, 4692, 4693, 4695: oled_data = 16'b0011101000001000;
         4713, 4720, 4722, 4723, 4725, 4730, 4731, 4733, 4734, 4735: oled_data = 16'b0011101000001000;
         4736, 4738, 4739, 4741, 4742, 4744, 4747, 4750, 4751, 4752: oled_data = 16'b0011101000001000;
         4754, 4758, 4763, 4765, 4768, 4769, 4771, 4772, 4774, 4776: oled_data = 16'b0011101000001000;
         4777, 4779, 4781, 4784, 4787, 4789, 4809, 4810, 4812, 4813: oled_data = 16'b0011101000001000;
         4814, 4880, 4882, 4883, 4885, 4907, 4910, 4977, 4980, 4982: oled_data = 16'b0011101000001000;
         4983, 5001, 5002, 5004, 5005, 5007, 5073, 5074, 5076, 5079: oled_data = 16'b0011101000001000;
         5097, 5099, 5102, 5169, 5173, 5174, 5193, 5194, 5195, 5199: oled_data = 16'b0011101000001000;
         5265, 5266, 5267, 5268, 5271, 5289, 5293, 5295, 5296, 5361: oled_data = 16'b0011101000001000;
         5365, 5366, 5386, 5388, 5390, 5392, 5457, 5458, 5460, 5461: oled_data = 16'b0011101000001000;
         5463, 5482, 5485, 5488, 5553, 5559, 5577, 5579, 5583, 5649: oled_data = 16'b0011101000001000;
         5650, 5652, 5653, 5655, 5676, 5679, 5680, 5745, 5749, 5769: oled_data = 16'b0011101000001000;
         5771, 5841, 5842, 5843, 5844, 5846, 5847, 5865, 5868, 5871: oled_data = 16'b0011101000001000;
         5872, 5937, 5941, 5966, 5968, 6033, 6035, 6037, 6057, 6059: oled_data = 16'b0011101000001000;
         6062, 6063, 6129, 6132, 6134, 6135: oled_data = 16'b0011101000001000;
         1939, 2031, 2122, 2135, 2198, 2379, 2390, 2582, 2806, 2996: oled_data = 16'b0111001111010001;
         3090, 3093, 3100, 3117, 5125, 5128: oled_data = 16'b0111001111010001;
         2008, 2096, 2392, 2488, 2776, 2872, 3064: oled_data = 16'b0110001101001110;
         2021, 5765: oled_data = 16'b1100111001111010;
         2032, 2095, 2613, 2968: oled_data = 16'b0110101110001110;
         2033, 2388, 2676: oled_data = 16'b0110001101001101;
         2040, 2087: oled_data = 16'b0111101110001110;
         2041, 2043, 2045, 2047, 2049, 2051, 2053, 2054, 2055, 2059: oled_data = 16'b0111101101001110;
         2060, 2062, 2064, 2066, 2068, 2069, 2071, 2073, 2074, 2076: oled_data = 16'b0111101101001110;
         2078, 2079, 2081, 2083, 2085, 2086: oled_data = 16'b0111101101001110;
         2042, 2044, 2046, 2048, 2050, 2052, 2056, 2058, 2061, 2063: oled_data = 16'b0111101101001101;
         2065, 2067, 2070, 2072, 2075, 2077, 2080, 2082, 2084: oled_data = 16'b0111101101001101;
         2057: oled_data = 16'b0111001101001110;
         2104, 2296, 2584, 2680, 3160: oled_data = 16'b0110101101001110;
         2120, 2228, 2416, 2479, 2513, 2576, 2708, 3080, 3484, 3486: oled_data = 16'b0011100111001000;
         3504, 3514, 3517, 3520, 3523, 3529, 3542, 3562, 3565, 3568: oled_data = 16'b0011100111001000;
         3570, 3572, 3574, 3576, 3577, 3579, 3581, 3583, 3587, 3589: oled_data = 16'b0011100111001000;
         3593, 3595, 3597, 3599, 3601, 3603, 3605, 3607, 3610, 3612: oled_data = 16'b0011100111001000;
         3616, 3618, 3620, 3622, 3624, 3626, 3628, 3632, 3634, 3635: oled_data = 16'b0011100111001000;
         3638, 3662, 3666, 3668, 3671, 3673, 3675, 3677, 3680, 3682: oled_data = 16'b0011100111001000;
         3685, 3688, 3691, 3693, 3695, 3697, 3699, 3701, 3703, 3705: oled_data = 16'b0011100111001000;
         3708, 3711, 3714, 3716, 3717, 3720, 3723, 3731, 3755, 3756: oled_data = 16'b0011100111001000;
         3852, 3926, 4042, 4044, 4047, 4052, 4058, 4075, 4083, 4093: oled_data = 16'b0011100111001000;
         4109, 4112, 4116, 4118, 4139, 4142, 4146, 4149, 4153, 4160: oled_data = 16'b0011100111001000;
         4162, 4169, 4177, 4180, 4182, 4193, 4195, 4199, 4201, 4236: oled_data = 16'b0011100111001000;
         4239, 4243, 4253, 4257, 4265, 4267, 4270, 4274, 4285, 4288: oled_data = 16'b0011100111001000;
         4303, 4306, 4330, 4333, 4343, 4345, 4350, 4352, 4355, 4359: oled_data = 16'b0011100111001000;
         4362, 4368, 4371, 4373, 4376, 4379, 4382, 4385, 4387, 4393: oled_data = 16'b0011100111001000;
         4395, 4400, 4403, 4430, 4436, 4440, 4444, 4449, 4459, 4462: oled_data = 16'b0011100111001000;
         4468, 4471, 4474, 4476, 4479, 4482, 4485, 4490, 4494, 4497: oled_data = 16'b0011100111001000;
         4500, 4524, 4530, 4533, 4535, 4538, 4543, 4546, 4553, 4556: oled_data = 16'b0011100111001000;
         4559, 4562, 4568, 4573, 4576, 4584, 4587, 4589, 4597, 4621: oled_data = 16'b0011100111001000;
         4624, 4632, 4640, 4646, 4648, 4654, 4659, 4665, 4667, 4669: oled_data = 16'b0011100111001000;
         4676, 4678, 4689, 4694, 4714, 4716, 4726, 4729, 4745, 4748: oled_data = 16'b0011100111001000;
         4756, 4759, 4783, 4791, 4815, 4884, 4886, 4906, 4912, 4976: oled_data = 16'b0011100111001000;
         4978, 5075, 5100, 5103, 5175, 5176, 5197, 5290, 5292, 5387: oled_data = 16'b0011100111001000;
         5459, 5481, 5486, 5557, 5578, 5581, 5651, 5675, 5678, 5773: oled_data = 16'b0011100111001000;
         5867, 5870, 5940, 5962, 5964, 6034, 6039, 6064, 6131: oled_data = 16'b0011100111001000;
         2126, 2189, 2701, 2896, 2959: oled_data = 16'b0101101100001100;
         2131, 5357, 5549, 5741, 5933, 6125: oled_data = 16'b0100001001001001;
         2136, 2232, 2279, 2328, 2471, 2520, 2616, 2663, 2759: oled_data = 16'b1010101000001000;
         2137, 2138, 2140, 2141, 2142, 2145, 2146, 2150, 2152, 2153: oled_data = 16'b1101000111000111;
         2154, 2156, 2157, 2158, 2159, 2161, 2162, 2163, 2165, 2166: oled_data = 16'b1101000111000111;
         2169, 2171, 2172, 2175, 2176, 2179, 2180, 2182, 2235, 2237: oled_data = 16'b1101000111000111;
         2239, 2240, 2243, 2244, 2245, 2246, 2252, 2257, 2259, 2263: oled_data = 16'b1101000111000111;
         2265, 2266, 2268, 2270, 2271, 2273, 2274, 2277, 2329, 2331: oled_data = 16'b1101000111000111;
         2332, 2333, 2334, 2336, 2337, 2339, 2341, 2343, 2344, 2345: oled_data = 16'b1101000111000111;
         2346, 2348, 2349, 2351, 2352, 2354, 2356, 2357, 2359, 2360: oled_data = 16'b1101000111000111;
         2362, 2363, 2364, 2365, 2367, 2368, 2370, 2371, 2373, 2425: oled_data = 16'b1101000111000111;
         2426, 2428, 2430, 2433, 2434, 2438, 2440, 2442, 2443, 2445: oled_data = 16'b1101000111000111;
         2446, 2447, 2449, 2450, 2451, 2453, 2454, 2456, 2457, 2458: oled_data = 16'b1101000111000111;
         2460, 2462, 2463, 2465, 2468, 2469, 2522, 2524, 2527, 2528: oled_data = 16'b1101000111000111;
         2530, 2532, 2533, 2536, 2537, 2539, 2540, 2545, 2547, 2550: oled_data = 16'b1101000111000111;
         2551, 2552, 2554, 2557, 2560, 2561, 2563, 2566, 2617, 2618: oled_data = 16'b1101000111000111;
         2620, 2622, 2623, 2625, 2626, 2627, 2629, 2630, 2632, 2634: oled_data = 16'b1101000111000111;
         2637, 2638, 2639, 2640, 2642, 2643, 2645, 2648, 2651, 2652: oled_data = 16'b1101000111000111;
         2653, 2655, 2657, 2658, 2660, 2661, 2662, 2713, 2715, 2716: oled_data = 16'b1101000111000111;
         2717, 2719, 2720, 2721, 2723, 2724, 2726, 2727, 2729, 2731: oled_data = 16'b1101000111000111;
         2732, 2733, 2737, 2738, 2741, 2743, 2744, 2746, 2747, 2749: oled_data = 16'b1101000111000111;
         2750, 2752, 2755: oled_data = 16'b1101000111000111;
         2139, 2143, 2147, 2149, 2151, 2155, 2160, 2164, 2167, 2170: oled_data = 16'b1101000111000110;
         2174, 2177, 2181, 2233, 2241, 2248, 2250, 2253, 2255, 2261: oled_data = 16'b1101000111000110;
         2264, 2269, 2275, 2278, 2330, 2335, 2338, 2340, 2342, 2347: oled_data = 16'b1101000111000110;
         2350, 2353, 2355, 2358, 2369, 2372, 2427, 2429, 2432, 2436: oled_data = 16'b1101000111000110;
         2439, 2448, 2452, 2459, 2461, 2464, 2467, 2470, 2521, 2526: oled_data = 16'b1101000111000110;
         2531, 2534, 2538, 2541, 2543, 2549, 2553, 2556, 2559, 2562: oled_data = 16'b1101000111000110;
         2565, 2619, 2621, 2624, 2628, 2631, 2633, 2636, 2641, 2644: oled_data = 16'b1101000111000110;
         2647, 2650, 2654, 2659, 2730, 2734, 2736, 2739, 2742, 2745: oled_data = 16'b1101000111000110;
         2751, 2753, 2756, 2758: oled_data = 16'b1101000111000110;
         2144, 2148, 2168, 2173, 2178, 2234, 2242, 2247, 2249, 2251: oled_data = 16'b1101001000000111;
         2254, 2256, 2260, 2262, 2276, 2374, 2431, 2435, 2437, 2466: oled_data = 16'b1101001000000111;
         2523, 2525, 2535, 2542, 2544, 2548, 2555, 2558, 2564, 2635: oled_data = 16'b1101001000000111;
         2646, 2649, 2656, 2728, 2735, 2740, 2754, 2757: oled_data = 16'b1101001000000111;
         2183, 2375, 2424, 2567, 2712: oled_data = 16'b1010001000001000;
         2203, 2299, 3163, 3259, 3835, 4027, 4699, 5275, 5467, 6139: oled_data = 16'b0111001100001101;
         2221, 2897, 2960: oled_data = 16'b0101101011001100;
         2236, 2238, 2258, 2267, 2272, 2361, 2366, 2441, 2444, 2455: oled_data = 16'b1101001000000110;
         2529, 2546, 2714, 2718, 2722, 2725, 2748: oled_data = 16'b1101001000000110;
         2284: oled_data = 16'b0110001100001101;
         2291, 3544, 3640, 3828, 4408, 5168, 5264, 5272, 5360, 5456: oled_data = 16'b0011000110000111;
         5552, 5648, 5744, 5840, 5936, 6032, 6136: oled_data = 16'b0011000110000111;
         2309, 2405, 2885, 3077, 3653, 3941, 4421, 4517, 4709, 5285: oled_data = 16'b1100110111111000;
         5381, 5957: oled_data = 16'b1100110111111000;
         2320, 2415: oled_data = 16'b0001000011000010;
         2325, 2412, 2898, 2961: oled_data = 16'b0110101110001111;
         2380, 2481, 2668, 3177, 3178, 3179, 3180, 3181, 3182, 3183: oled_data = 16'b0010100101000101;
         3184, 3185, 3186, 3187, 3189, 3190, 3191, 3192, 3193, 3194: oled_data = 16'b0010100101000101;
         3195, 3196, 3197, 3198, 3199, 3201, 3202, 3203, 3204, 3206: oled_data = 16'b0010100101000101;
         3207, 3208, 3209, 3210, 3211, 3212, 3214, 3215, 3217, 3218: oled_data = 16'b0010100101000101;
         3220, 3221, 3222, 3223, 3224, 3225, 3226, 3227, 3228, 3229: oled_data = 16'b0010100101000101;
         3230, 3231, 3232, 3233, 3234, 3235, 3236, 3238, 3239, 3240: oled_data = 16'b0010100101000101;
         3241, 3242, 3244, 3246, 3247, 3248, 3249, 3251, 3252, 3253: oled_data = 16'b0010100101000101;
         3254, 3255, 3924: oled_data = 16'b0010100101000101;
         2383, 5105, 5393, 5873: oled_data = 16'b0001100010000011;
         2408, 2792, 3658, 3829, 3850, 4145, 4151, 4158, 4164, 4167: oled_data = 16'b0100000111001000;
         4172, 4184, 4186, 4191, 4197, 4203, 4206, 4209, 4278, 4309: oled_data = 16'b0100000111001000;
         4338, 4341, 4347, 4522, 4579, 4592, 4595, 4638, 4686, 4718: oled_data = 16'b0100000111001000;
         4721, 4724, 4737, 4773, 4775, 5294, 5484, 5942, 6061, 6133: oled_data = 16'b0100000111001000;
         2417, 3561, 3571, 3578, 3588, 3598, 3602, 3606, 3611, 3617: oled_data = 16'b0011101000001001;
         3633, 3659, 3830, 3849, 3851, 4021, 4046, 4049, 4051, 4053: oled_data = 16'b0011101000001001;
         4055, 4057, 4059, 4062, 4064, 4066, 4068, 4072, 4074, 4076: oled_data = 16'b0011101000001001;
         4081, 4084, 4087, 4089, 4091, 4094, 4097, 4099, 4101, 4104: oled_data = 16'b0011101000001001;
         4106, 4108, 4110, 4113, 4141, 4144, 4178, 4181, 4192, 4198: oled_data = 16'b0011101000001001;
         4207, 4213, 4235, 4242, 4244, 4248, 4254, 4256, 4258, 4264: oled_data = 16'b0011101000001001;
         4266, 4268, 4272, 4279, 4286, 4290, 4298, 4305, 4332, 4334: oled_data = 16'b0011101000001001;
         4348, 4370, 4372, 4374, 4378, 4384, 4404, 4425, 4435, 4437: oled_data = 16'b0011101000001001;
         4439, 4441, 4443, 4446, 4448, 4450, 4458, 4460, 4463, 4472: oled_data = 16'b0011101000001001;
         4477, 4481, 4483, 4489, 4491, 4496, 4558, 4563, 4569, 4580: oled_data = 16'b0011101000001001;
         4590, 4594, 4596, 4598, 4617, 4619, 4625, 4629, 4631, 4633: oled_data = 16'b0011101000001001;
         4639, 4641, 4647, 4649, 4653, 4677, 4679, 4688, 4717, 4719: oled_data = 16'b0011101000001001;
         4728, 4755, 4757, 4760, 4782, 4816, 4887, 5008, 5196, 5198: oled_data = 16'b0011101000001001;
         5389, 5483, 5556, 5580, 5582, 5673, 5772, 5774, 5943, 5961: oled_data = 16'b0011101000001001;
         5963, 5965, 6036, 6038, 6060: oled_data = 16'b0011101000001001;
         2421: oled_data = 16'b0101001010001010;
         2484, 5453, 5837: oled_data = 16'b0100101001001001;
         2508: oled_data = 16'b0111001111001111;
         2511: oled_data = 16'b0001100010000010;
         2514, 3656, 3752, 3944, 4040, 4232, 4520, 4712, 4808, 5096: oled_data = 16'b0010000100000101;
         5192, 5288, 5864: oled_data = 16'b0010000100000101;
         2517: oled_data = 16'b0100101010001010;
         2577, 3256, 5480: oled_data = 16'b0010000101000101;
         2580: oled_data = 16'b0100101001001010;
         2597, 3269, 5573: oled_data = 16'b1100111001111001;
         2764: oled_data = 16'b0101101100001101;
         2771, 5072, 6128: oled_data = 16'b0011000110000110;
         2798: oled_data = 16'b0101001011001011;
         2803, 3467, 3470, 3473, 3476, 3478, 3480, 3482, 3489, 3492: oled_data = 16'b0011100111000111;
         3495, 3498, 3500, 3502, 3506, 3508, 3510, 3526, 3532, 3535: oled_data = 16'b0011100111000111;
         3538, 3540, 3663, 3665, 3669, 3679, 3683, 3686, 3689, 3707: oled_data = 16'b0011100111000111;
         3710, 3713, 3719, 3722, 3725, 3726, 3728, 3729, 4020, 4216: oled_data = 16'b0011100111000111;
         4792, 5165, 5368, 6040: oled_data = 16'b0011100111000111;
         2808, 2855: oled_data = 16'b1001001010001010;
         2809, 2812, 2814, 2815, 2817, 2818, 2819, 2821, 2822, 2825: oled_data = 16'b1010001001001001;
         2826, 2828, 2830, 2832, 2834, 2836, 2837, 2839, 2842, 2843: oled_data = 16'b1010001001001001;
         2846, 2847, 2849, 2851, 2853, 2854: oled_data = 16'b1010001001001001;
         2810, 2813, 2820, 2824, 2829, 2831, 2833, 2835, 2838, 2841: oled_data = 16'b1010101001001001;
         2844, 2848, 2852: oled_data = 16'b1010101001001001;
         2811, 2823, 2840, 2845, 2850: oled_data = 16'b1010001001001000;
         2816, 2827: oled_data = 16'b1010101001001000;
         2861: oled_data = 16'b0101001011001100;
         2866, 3465, 3468, 3471, 3475, 3483, 3485, 3487, 3490, 3493: oled_data = 16'b0011000111000111;
         3496, 3503, 3505, 3511, 3513, 3515, 3516, 3518, 3519, 3521: oled_data = 16'b0011000111000111;
         3522, 3524, 3528, 3530, 3534, 3537, 3541, 3543, 3667, 3672: oled_data = 16'b0011000111000111;
         3674, 3676, 3681, 3684, 3687, 3692, 3694, 3696, 3698, 3700: oled_data = 16'b0011000111000111;
         3702, 3704, 3706, 3709, 3712, 3715, 3736, 3832, 4024, 4120: oled_data = 16'b0011000111000111;
         4312, 4504, 4696, 4817, 4888, 5080, 5464, 5656, 5752, 5944: oled_data = 16'b0011000111000111;
         3188, 3200, 3205, 3216, 3219, 3237, 3243, 3250, 4879: oled_data = 16'b0010100101000110;
         3213, 3245: oled_data = 16'b0010100110000101;
         3466, 3469, 3472, 3474, 3477, 3479, 3481, 3488, 3491, 3494: oled_data = 16'b0011000111001000;
         3497, 3499, 3501, 3507, 3509, 3525, 3527, 3531, 3533, 3536: oled_data = 16'b0011000111001000;
         3539, 3664, 3670, 3678, 3690, 3718, 3721, 3724, 3727, 3730: oled_data = 16'b0011000111001000;
         3512: oled_data = 16'b0011100110001000;
         3557, 4997: oled_data = 16'b1101011001111010;
         3564, 3567, 3585, 3591, 3614, 3630, 3637, 4023, 4070, 4078: oled_data = 16'b0011100111001001;
         4175, 4215, 4246, 4250, 4260, 4262, 4281, 4292, 4296, 4300: oled_data = 16'b0011100111001001;
         4336, 4365, 4390, 4406, 4427, 4433, 4452, 4454, 4456, 4465: oled_data = 16'b0011100111001001;
         4487, 4503, 4527, 4541, 4549, 4565, 4627, 4643, 4651, 4656: oled_data = 16'b0011100111001001;
         4662, 4671, 4673, 4681, 4732, 4753, 4762, 4766, 4780, 4786: oled_data = 16'b0011100111001001;
         4811, 4881, 4909, 4981, 5003, 5006, 5078, 5170, 5172, 5200: oled_data = 16'b0011100111001001;
         5269, 5362, 5364, 5367, 5391, 5462, 5554, 5584, 5654, 5746: oled_data = 16'b0011100111001001;
         5748, 5751, 5770, 5776, 5845, 5938, 5967: oled_data = 16'b0011100111001001;
         3735, 4137, 4156, 4188, 4211, 4397, 4635, 4740, 4770, 4778: oled_data = 16'b0100000111001001;
         4788, 5098: oled_data = 16'b0100000111001001;
         3749: oled_data = 16'b1100110110111000;
         3928, 4600, 4984, 5560, 5848: oled_data = 16'b0011100110000111;
         3949: oled_data = 16'b0010100100000101;
         4043, 4380, 4399, 4402, 4525, 4571, 4574, 4588, 4746, 4764: oled_data = 16'b0100001000001001;
         4790, 4905, 4979, 5261, 5291, 5385, 5645, 6029, 6130: oled_data = 16'b0100001000001001;
         4136: oled_data = 16'b0010000101000100;
         5201, 5585, 5777: oled_data = 16'b0001100011000010;
         5204, 5396, 5588, 5780, 5972: oled_data = 16'b1001110011110101;
         5205, 5207, 5209, 5211, 5213, 5215, 5217, 5219, 5221, 5223: oled_data = 16'b1001110100110101;
         5225, 5227, 5229, 5231, 5233, 5235, 5237, 5239, 5241, 5243: oled_data = 16'b1001110100110101;
         5245, 5247, 5249, 5251, 5253, 5255, 5257, 5259, 5302, 5304: oled_data = 16'b1001110100110101;
         5306, 5308, 5310, 5312, 5318, 5320, 5324, 5326, 5328, 5330: oled_data = 16'b1001110100110101;
         5332, 5334, 5336, 5338, 5340, 5342, 5344, 5348, 5350, 5354: oled_data = 16'b1001110100110101;
         5356, 5397, 5399, 5403, 5405, 5407, 5409, 5411, 5413, 5415: oled_data = 16'b1001110100110101;
         5417, 5419, 5421, 5429, 5431, 5433, 5435, 5439, 5441, 5445: oled_data = 16'b1001110100110101;
         5447, 5449, 5451, 5493, 5495, 5497, 5501, 5503, 5505, 5511: oled_data = 16'b1001110100110101;
         5515, 5517, 5519, 5522, 5524, 5526, 5528, 5531, 5533, 5540: oled_data = 16'b1001110100110101;
         5548, 5594, 5596, 5598, 5604, 5606, 5608, 5610, 5612, 5623: oled_data = 16'b1001110100110101;
         5627, 5631, 5634, 5635, 5637, 5639, 5641, 5685, 5687, 5689: oled_data = 16'b1001110100110101;
         5691, 5695, 5697, 5699, 5707, 5709, 5711, 5713, 5715, 5717: oled_data = 16'b1001110100110101;
         5720, 5722, 5724, 5728, 5730, 5732, 5736, 5738, 5740, 5784: oled_data = 16'b1001110100110101;
         5786, 5791, 5794, 5796, 5798, 5800, 5802, 5804, 5812, 5814: oled_data = 16'b1001110100110101;
         5816, 5823, 5825, 5829, 5832, 5834, 5879, 5883, 5887, 5889: oled_data = 16'b1001110100110101;
         5891, 5893, 5896, 5901, 5903, 5905, 5907, 5909, 5911, 5913: oled_data = 16'b1001110100110101;
         5915, 5917, 5919, 5921, 5926, 5928, 5930, 5932, 5973, 5975: oled_data = 16'b1001110100110101;
         5977, 5980, 5982, 5988, 5990, 5992, 5994, 5998, 6001, 6007: oled_data = 16'b1001110100110101;
         6009, 6011, 6013, 6015, 6019, 6021, 6023, 6025, 6027, 6070: oled_data = 16'b1001110100110101;
         6072, 6074, 6076, 6078, 6080, 6082, 6084, 6086, 6088, 6090: oled_data = 16'b1001110100110101;
         6092, 6095, 6097, 6099, 6101, 6105, 6107, 6109, 6111, 6113: oled_data = 16'b1001110100110101;
         6115, 6117, 6121, 6123: oled_data = 16'b1001110100110101;
         5206, 5208, 5210, 5212, 5214, 5216, 5218, 5220, 5222, 5224: oled_data = 16'b1001110100110110;
         5226, 5228, 5230, 5232, 5234, 5236, 5238, 5240, 5242, 5244: oled_data = 16'b1001110100110110;
         5246, 5248, 5250, 5252, 5254, 5256, 5258, 5260, 5301, 5303: oled_data = 16'b1001110100110110;
         5305, 5307, 5309, 5311, 5313, 5315, 5321, 5323, 5327, 5329: oled_data = 16'b1001110100110110;
         5331, 5333, 5335, 5337, 5341, 5345, 5347, 5351, 5353, 5400: oled_data = 16'b1001110100110110;
         5402, 5410, 5412, 5414, 5416, 5418, 5422, 5424, 5426, 5428: oled_data = 16'b1001110100110110;
         5434, 5436, 5438, 5440, 5442, 5444, 5446, 5448, 5450, 5452: oled_data = 16'b1001110100110110;
         5494, 5496, 5498, 5502, 5504, 5506, 5508, 5510, 5516, 5518: oled_data = 16'b1001110100110110;
         5520, 5521, 5523, 5525, 5527, 5529, 5532, 5534, 5538, 5539: oled_data = 16'b1001110100110110;
         5543, 5547, 5589, 5591, 5593, 5595, 5597, 5601, 5603, 5605: oled_data = 16'b1001110100110110;
         5609, 5611, 5615, 5617, 5620, 5626, 5630, 5632, 5633, 5638: oled_data = 16'b1001110100110110;
         5640, 5642, 5643, 5686, 5688, 5692, 5694, 5696, 5698, 5702: oled_data = 16'b1001110100110110;
         5704, 5706, 5710, 5712, 5714, 5716, 5718, 5721, 5723, 5725: oled_data = 16'b1001110100110110;
         5727, 5731, 5733, 5735, 5739, 5781, 5785, 5787, 5789, 5790: oled_data = 16'b1001110100110110;
         5793, 5797, 5799, 5801, 5803, 5805, 5807, 5809, 5811, 5815: oled_data = 16'b1001110100110110;
         5817, 5819, 5821, 5822, 5824, 5826, 5828, 5830, 5831, 5833: oled_data = 16'b1001110100110110;
         5836, 5878, 5880, 5882, 5884, 5888, 5892, 5895, 5898, 5900: oled_data = 16'b1001110100110110;
         5902, 5904, 5906, 5908, 5910, 5914, 5916, 5922, 5924, 5931: oled_data = 16'b1001110100110110;
         5974, 5976, 5978, 5981, 5983, 5985, 5987, 5989, 5991, 5993: oled_data = 16'b1001110100110110;
         5995, 5999, 6002, 6006, 6008, 6014, 6016, 6020, 6022, 6024: oled_data = 16'b1001110100110110;
         6026, 6069, 6079, 6081, 6091, 6093, 6094, 6096, 6098, 6100: oled_data = 16'b1001110100110110;
         6102, 6106, 6112, 6114, 6118, 6120, 6124: oled_data = 16'b1001110100110110;
         5300, 5684: oled_data = 16'b1001010011110101;
         5314, 5322, 5346, 5352, 5401, 5423, 5425, 5427, 5437, 5443: oled_data = 16'b1010010100110101;
         5499, 5507, 5509, 5535, 5537, 5542, 5544, 5546, 5590, 5602: oled_data = 16'b1010010100110101;
         5616, 5621, 5644, 5693, 5701, 5703, 5705, 5726, 5734, 5788: oled_data = 16'b1010010100110101;
         5806, 5808, 5810, 5818, 5820, 5827, 5877, 5881, 5899, 5984: oled_data = 16'b1010010100110101;
         6003, 6005, 6103, 6119: oled_data = 16'b1010010100110101;
         5316, 5513, 5600, 5614, 5618, 5625, 5629, 5782, 5885, 5923: oled_data = 16'b1001110101110101;
         5986, 5996, 6017: oled_data = 16'b1001110101110101;
         5317, 5319, 5325, 5339, 5343, 5349, 5355, 5398, 5404, 5406: oled_data = 16'b1010010100110110;
         5408, 5420, 5430, 5432, 5512, 5514, 5530, 5599, 5613, 5619: oled_data = 16'b1010010100110110;
         5624, 5628, 5636, 5690, 5708, 5719, 5729, 5737, 5783, 5792: oled_data = 16'b1010010100110110;
         5795, 5813, 5835, 5886, 5890, 5894, 5897, 5912, 5918, 5920: oled_data = 16'b1010010100110110;
         5925, 5929, 5979, 5997, 6010, 6018, 6028, 6071, 6073, 6077: oled_data = 16'b1010010100110110;
         6083, 6085, 6087, 6089, 6108, 6110, 6116, 6122: oled_data = 16'b1010010100110110;
         5492, 5876, 6068: oled_data = 16'b1001010100110101;
         5500, 5536, 5541, 5545, 5607, 5622, 5700, 6004, 6012, 6075: oled_data = 16'b1001110101110110;
         6104: oled_data = 16'b1001110101110110;
         5592: oled_data = 16'b1010010101110101;
         5669: oled_data = 16'b1101011010111010;
         5927, 6000: oled_data = 16'b1010010101110110;
         6053: oled_data = 16'b1101010110111000;
         default: oled_data = 16'b0000000000000000;
     endcase end end endmodule
