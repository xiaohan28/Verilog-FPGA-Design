`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.10.2024 15:23:34
// Design Name: 
// Module Name: frame_data_feature2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tryagain( 
    output reg [15:0] oled_data,
    input frame_rate, 
    input [12:0] pixel_index  
    );
    

    // lives
    always @ (posedge frame_rate) begin
        case (pixel_index)
        0, 2, 5, 9, 12, 14, 15, 17, 20, 24: oled_data = 16'b1111111100111101;
        27, 29, 30, 32, 35, 39, 42, 44, 45, 47: oled_data = 16'b1111111100111101;
        50, 54, 57, 59, 60, 62, 65, 69, 72, 74: oled_data = 16'b1111111100111101;
        75, 77, 80, 84, 87, 89, 90, 92, 95, 96: oled_data = 16'b1111111100111101;
        99, 103, 106, 108, 109, 111, 114, 118, 121, 123: oled_data = 16'b1111111100111101;
        124, 126, 129, 133, 136, 138, 139, 141, 144, 148: oled_data = 16'b1111111100111101;
        151, 153, 154, 156, 159, 163, 166, 168, 169, 171: oled_data = 16'b1111111100111101;
        174, 178, 181, 183, 184, 186, 189, 194, 196, 197: oled_data = 16'b1111111100111101;
        199, 202, 206, 209, 211, 212, 214, 217, 221, 224: oled_data = 16'b1111111100111101;
        226, 227, 229, 232, 236, 239, 241, 242, 244, 247: oled_data = 16'b1111111100111101;
        251, 254, 256, 257, 259, 262, 266, 269, 271, 272: oled_data = 16'b1111111100111101;
        274, 277, 281, 284, 286, 288, 290, 291, 293, 299: oled_data = 16'b1111111100111101;
        301, 303, 309, 311, 313, 319, 321, 323, 329, 331: oled_data = 16'b1111111100111101;
        333, 339, 341, 343, 349, 351, 353, 359, 361, 363: oled_data = 16'b1111111100111101;
        369, 371, 373, 379, 381, 383, 384, 390, 393, 397: oled_data = 16'b1111111100111101;
        400, 402, 405, 408, 412, 417, 418, 420, 430, 432: oled_data = 16'b1111111100111101;
        433, 438, 442, 445, 448, 450, 453, 457, 460, 462: oled_data = 16'b1111111100111101;
        465, 468, 472, 477, 483, 487, 489, 491, 492, 494: oled_data = 16'b1111111100111101;
        497, 499, 502, 507, 511, 516, 519, 521, 524, 526: oled_data = 16'b1111111100111101;
        527, 529, 531, 532, 534, 537, 539, 542, 547, 551: oled_data = 16'b1111111100111101;
        556, 559, 561, 564, 566, 567, 569, 571, 572, 574: oled_data = 16'b1111111100111101;
        576, 578, 580, 581, 584, 593, 595, 600, 606, 608: oled_data = 16'b1111111100111101;
        611, 613, 615, 616, 618, 620, 625, 631, 636, 638: oled_data = 16'b1111111100111101;
        640, 641, 643, 645, 648, 650, 656, 661, 663, 666: oled_data = 16'b1111111100111101;
        668, 670, 675, 678, 681, 682, 685, 686, 689, 690: oled_data = 16'b1111111100111101;
        692, 694, 697, 699, 702, 705, 709, 710, 712, 714: oled_data = 16'b1111111100111101;
        715, 717, 719, 722, 724, 725, 729, 730, 734, 735: oled_data = 16'b1111111100111101;
        737, 740, 742, 744, 745, 747, 749, 750, 754, 757: oled_data = 16'b1111111100111101;
        760, 762, 765, 767, 768, 770, 772, 779, 787, 789: oled_data = 16'b1111111100111101;
        791, 793, 796, 798, 803, 809, 811, 814, 816, 818: oled_data = 16'b1111111100111101;
        819, 821, 823, 828, 834, 839, 841, 843, 844, 846: oled_data = 16'b1111111100111101;
        848, 851, 853, 859, 864, 867, 869, 871, 874, 877: oled_data = 16'b1111111100111101;
        880, 883, 886, 895, 897, 900, 903, 907, 912, 913: oled_data = 16'b1111111100111101;
        915, 918, 925, 927, 928, 937, 943, 945, 948, 955: oled_data = 16'b1111111100111101;
        957, 962, 964, 969, 971, 974, 976, 980, 983, 986: oled_data = 16'b1111111100111101;
        988, 990, 997, 999, 1002, 1004, 1006, 1007, 1009, 1011: oled_data = 16'b1111111100111101;
        1016, 1019, 1022, 1027, 1029, 1031, 1032, 1034, 1036, 1039: oled_data = 16'b1111111100111101;
        1041, 1047, 1051, 1052, 1054, 1055, 1056, 1058, 1059, 1062: oled_data = 16'b1111111100111101;
        1065, 1067, 1071, 1073, 1075, 1077, 1080, 1083, 1085, 1086: oled_data = 16'b1111111100111101;
        1088, 1089, 1091, 1093, 1096, 1101, 1105, 1108, 1110, 1113: oled_data = 16'b1111111100111101;
        1115, 1118, 1120, 1121, 1123, 1125, 1126, 1128, 1131, 1133: oled_data = 16'b1111111100111101;
        1136, 1140, 1141, 1145, 1150, 1152, 1162, 1179, 1183, 1185: oled_data = 16'b1111111100111101;
        1186, 1188, 1195, 1199, 1202, 1204, 1210, 1212, 1214, 1215: oled_data = 16'b1111111100111101;
        1217, 1220, 1222, 1224, 1227, 1230, 1234, 1240, 1242, 1244: oled_data = 16'b1111111100111101;
        1247, 1251, 1253, 1256, 1258, 1261, 1275, 1277, 1280, 1282: oled_data = 16'b1111111100111101;
        1283, 1285, 1286, 1289, 1292, 1294, 1296, 1298, 1299, 1301: oled_data = 16'b1111111100111101;
        1303, 1306, 1308, 1314, 1318, 1319, 1321, 1324, 1326, 1328: oled_data = 16'b1111111100111101;
        1331, 1333, 1334, 1344, 1346, 1348, 1350, 1352, 1353, 1355: oled_data = 16'b1111111100111101;
        1425, 1427, 1428, 1430, 1437, 1448, 1451, 1521, 1527, 1529: oled_data = 16'b1111111100111101;
        1531, 1534, 1536, 1538, 1540, 1543, 1546, 1548, 1617, 1620: oled_data = 16'b1111111100111101;
        1621, 1623, 1626, 1628, 1630, 1632, 1635, 1637, 1638, 1640: oled_data = 16'b1111111100111101;
        1642, 1643, 1718, 1720, 1724, 1726, 1730, 1732, 1736, 1737: oled_data = 16'b1111111100111101;
        1739, 1740, 1810, 1811, 1813, 1815, 1817, 1820, 1824, 1826: oled_data = 16'b1111111100111101;
        1827, 1829, 1908, 1910, 1913, 1919, 1920, 1927, 1929, 1930: oled_data = 16'b1111111100111101;
        1932, 1933, 2002, 2004, 2008, 2010, 2013, 2019, 2021, 2024: oled_data = 16'b1111111100111101;
        2028, 2030, 2032, 2097, 2099, 2102, 2104, 2107, 2110, 2112: oled_data = 16'b1111111100111101;
        2114, 2116, 2119, 2121, 2124, 2126, 2129, 2192, 2195, 2197: oled_data = 16'b1111111100111101;
        2199, 2201, 2203, 2207, 2213, 2219, 2221, 2223, 2224, 2289: oled_data = 16'b1111111100111101;
        2291, 2294, 2300, 2301, 2303, 2304, 2306, 2310, 2312, 2315: oled_data = 16'b1111111100111101;
        2317, 2320, 2322, 2326, 2329, 2331, 2335, 2338, 2342, 2346: oled_data = 16'b1111111100111101;
        2348, 2358, 2360, 2366, 2368, 2376, 2378, 2382, 2389, 2391: oled_data = 16'b1111111100111101;
        2394, 2400, 2403, 2405, 2409, 2411, 2415, 2419, 2421, 2423: oled_data = 16'b1111111100111101;
        2426, 2428, 2432, 2437, 2440, 2443, 2445, 2449, 2450, 2452: oled_data = 16'b1111111100111101;
        2455, 2457, 2460, 2466, 2468, 2469, 2473, 2475, 2479, 2483: oled_data = 16'b1111111100111101;
        2486, 2488, 2491, 2493, 2498, 2500, 2502, 2505, 2509, 2511: oled_data = 16'b1111111100111101;
        2512, 2514, 2515, 2518, 2521, 2523, 2526, 2529, 2532, 2534: oled_data = 16'b1111111100111101;
        2537, 2539, 2543, 2544, 2546, 2548, 2550, 2554, 2557, 2560: oled_data = 16'b1111111100111101;
        2562, 2563, 2565, 2567, 2570, 2573, 2577, 2579, 2582, 2585: oled_data = 16'b1111111100111101;
        2587, 2588, 2591, 2592, 2594, 2597, 2599, 2605, 2609, 2611: oled_data = 16'b1111111100111101;
        2615, 2618, 2621, 2623, 2626, 2629, 2631, 2633, 2636, 2639: oled_data = 16'b1111111100111101;
        2641, 2643, 2644, 2646, 2648, 2650, 2652, 2654, 2656, 2657: oled_data = 16'b1111111100111101;
        2659, 2662, 2664, 2668, 2670, 2672, 2674, 2677, 2679, 2683: oled_data = 16'b1111111100111101;
        2685, 2688, 2692, 2696, 2698, 2700, 2702, 2703, 2705, 2706: oled_data = 16'b1111111100111101;
        2708, 2709, 2711, 2718, 2725, 2727, 2730, 2732, 2736, 2743: oled_data = 16'b1111111100111101;
        2746, 2747, 2749, 2758, 2760, 2762, 2766, 2769, 2771, 2775: oled_data = 16'b1111111100111101;
        2777, 2778, 2782, 2786, 2789, 2790, 2794, 2795, 2797, 2799: oled_data = 16'b1111111100111101;
        2810, 2816, 2819, 2824, 2827, 2829, 2830, 2840, 2846, 2859: oled_data = 16'b1111111100111101;
        2864, 2868, 2871, 2872, 2877, 2879, 2880, 2882, 2884, 2893: oled_data = 16'b1111111100111101;
        2896, 2913, 2921, 2923, 2924, 2926, 2927, 2931, 2935, 2942: oled_data = 16'b1111111100111101;
        2956, 2958, 2961, 2965, 2967, 2969, 2971, 2975, 2976, 2978: oled_data = 16'b1111111100111101;
        2979, 2981, 2985, 2987, 2988, 2990, 2992, 3018, 3020, 3027: oled_data = 16'b1111111100111101;
        3031, 3039, 3052, 3055, 3058, 3061, 3064, 3066, 3068, 3072: oled_data = 16'b1111111100111101;
        3076, 3078, 3081, 3090, 3096, 3097, 3102, 3114, 3115, 3117: oled_data = 16'b1111111100111101;
        3119, 3123, 3135, 3137, 3141, 3147, 3149, 3155, 3159, 3161: oled_data = 16'b1111111100111101;
        3163, 3165, 3166, 3170, 3175, 3178, 3181, 3182, 3186, 3210: oled_data = 16'b1111111100111101;
        3212, 3213, 3223, 3227, 3232, 3238, 3239, 3246, 3249, 3254: oled_data = 16'b1111111100111101;
        
        3256, 3257, 3259, 3260, 3263, 3264, 3266, 3269, 3280, 3302: oled_data = 16'b1111111100111101;
        3306, 3311, 3323, 3328, 3329, 3333, 3335, 3339, 3343, 3347: oled_data = 16'b1111111100111101;
        3351, 3353, 3354, 3356, 3357, 3360, 3363, 3365, 3367, 3368: oled_data = 16'b1111111100111101;
        3371, 3374, 3378, 3384, 3385, 3398, 3402, 3405, 3423, 3425: oled_data = 16'b1111111100111101;
        3436, 3437, 3439, 3445, 3448, 3450, 3465, 3467, 3471, 3474: oled_data = 16'b1111111100111101;
        3499, 3503, 3507, 3511, 3519, 3520, 3525, 3534, 3536, 3537: oled_data = 16'b1111111100111101;
        3540, 3542, 3545, 3550, 3552, 3554, 3557, 3558, 3561, 3565: oled_data = 16'b1111111100111101;
        3568, 3570, 3576, 3586, 3598, 3603, 3622, 3623, 3629, 3631: oled_data = 16'b1111111100111101;
        3633, 3636, 3638, 3643, 3647, 3660, 3662, 3663, 3665, 3667: oled_data = 16'b1111111100111101;
        3673, 3674, 3676, 3680, 3689, 3691, 3692, 3695, 3700, 3703: oled_data = 16'b1111111100111101;
        3712, 3717, 3719, 3723, 3726, 3730, 3732, 3735, 3736, 3738: oled_data = 16'b1111111100111101;
        3741, 3743, 3744, 3746, 3751, 3754, 3758, 3761, 3764, 3766: oled_data = 16'b1111111100111101;
        3768, 3770, 3771, 3773, 3775, 3777, 3778, 3781, 3783, 3784: oled_data = 16'b1111111100111101;
        3792, 3793, 3795, 3796, 3797, 3799, 3801, 3803, 3805, 3809: oled_data = 16'b1111111100111101;
        3815, 3821, 3824, 3826, 3827, 3833, 3835, 3837, 3840, 3845: oled_data = 16'b1111111100111101;
        3848, 3854, 3855, 3858, 3861, 3863, 3868, 3870, 3872, 3874: oled_data = 16'b1111111100111101;
        3878, 3881, 3883, 3887, 3889, 3895, 3896, 3898, 3899, 3900: oled_data = 16'b1111111100111101;
        3902, 3903, 3905, 3908, 3910, 3912, 3913, 3915, 3918, 3920: oled_data = 16'b1111111100111101;
        3921, 3926, 3929, 3930, 3932, 3934, 3935, 3938, 3942, 3944: oled_data = 16'b1111111100111101;
        3948, 3950, 3952, 3953, 3955, 3957, 3960, 3962, 3965, 3967: oled_data = 16'b1111111100111101;
        3969, 3973, 3975, 3977, 3978, 3980, 3982, 3984, 3986, 3987: oled_data = 16'b1111111100111101;
        3989, 3997, 3999, 4000, 4002, 4005, 4007, 4009, 4010, 4012: oled_data = 16'b1111111100111101;
        4015, 4017, 4019, 4023, 4028, 4032, 4034, 4037, 4039, 4042: oled_data = 16'b1111111100111101;
        4045, 4049, 4051, 4054, 4056, 4057, 4059, 4062, 4064, 4066: oled_data = 16'b1111111100111101;
        4070, 4072, 4074, 4077, 4079, 4080, 4084, 4088, 4090, 4092: oled_data = 16'b1111111100111101;
        4098, 4100, 4109, 4113, 4117, 4123, 4125, 4128, 4131, 4134: oled_data = 16'b1111111100111101;
        4136, 4138, 4140, 4156, 4160, 4162, 4165, 4167, 4171, 4177: oled_data = 16'b1111111100111101;
        4187, 4195, 4203, 4210, 4213, 4215, 4216, 4219, 4222, 4233: oled_data = 16'b1111111100111101;
        4235, 4257, 4262, 4264, 4266, 4268, 4274, 4283, 4284, 4290: oled_data = 16'b1111111100111101;
        4295, 4308, 4310, 4312, 4316, 4318, 4320, 4322, 4325, 4326: oled_data = 16'b1111111100111101;
        4330, 4332, 4359, 4371, 4387, 4401, 4404, 4406, 4409, 4413: oled_data = 16'b1111111100111101;
        4415, 4420, 4422, 4423, 4427, 4429, 4458, 4471, 4475, 4479: oled_data = 16'b1111111100111101;
        4487, 4498, 4503, 4505, 4506, 4508, 4510, 4512, 4514, 4520: oled_data = 16'b1111111100111101;
        4524, 4550, 4551, 4555, 4563, 4579, 4593, 4595, 4597, 4599: oled_data = 16'b1111111100111101;
        4600, 4602, 4605, 4607, 4608, 4610, 4613, 4618, 4621, 4644: oled_data = 16'b1111111100111101;
        4646, 4648, 4667, 4675, 4679, 4692, 4694, 4696, 4698, 4702: oled_data = 16'b1111111100111101;
        4707, 4714, 4742, 4746, 4771, 4779, 4786, 4789, 4797, 4799: oled_data = 16'b1111111100111101;
        4800, 4802, 4808, 4812, 4814, 4839, 4842, 4843, 4859, 4867: oled_data = 16'b1111111100111101;
        4871, 4876, 4882, 4886, 4889, 4891, 4892, 4894, 4896, 4899: oled_data = 16'b1111111100111101;
        4901, 4902, 4904, 4908, 4909, 4937, 4939, 4948, 4971, 4972: oled_data = 16'b1111111100111101;
        4979, 4980, 4986, 4988, 4989, 4991, 4994, 4996, 4998, 5002: oled_data = 16'b1111111100111101;
        
        5004, 5006, 5011, 5013, 5017, 5030, 5031, 5033, 5036, 5050: oled_data = 16'b1111111100111101;
        5052, 5056, 5059, 5060, 5064, 5073, 5078, 5080, 5082, 5086: oled_data = 16'b1111111100111101;
        5088, 5090, 5095, 5098, 5101, 5103, 5105, 5106, 5108, 5110: oled_data = 16'b1111111100111101;
        5118, 5124, 5125, 5127, 5128, 5130, 5132, 5135, 5136, 5138: oled_data = 16'b1111111100111101;
        5142, 5144, 5147, 5152, 5154, 5156, 5158, 5161, 5162, 5164: oled_data = 16'b1111111100111101;
        5166, 5168, 5170, 5174, 5177, 5179, 5181, 5183, 5184, 5186: oled_data = 16'b1111111100111101;
        5188, 5189, 5203, 5207, 5210, 5213, 5215, 5217, 5219, 5226: oled_data = 16'b1111111100111101;
        5229, 5233, 5235, 5236, 5238, 5239, 5241, 5245, 5249, 5252: oled_data = 16'b1111111100111101;
        5255, 5256, 5258, 5263, 5267, 5268, 5270, 5272, 5274, 5278: oled_data = 16'b1111111100111101;
        5280, 5283, 5286, 5288, 5289, 5291, 5292, 5295, 5297, 5300: oled_data = 16'b1111111100111101;
        5304, 5307, 5310, 5312, 5314, 5318, 5322, 5327, 5330, 5332: oled_data = 16'b1111111100111101;
        5333, 5335, 5336, 5338, 5339, 5341, 5344, 5346, 5352, 5355: oled_data = 16'b1111111100111101;
        5357, 5359, 5365, 5367, 5368, 5375, 5378, 5380, 5382, 5386: oled_data = 16'b1111111100111101;
        5388, 5391, 5398, 5402, 5404, 5406, 5409, 5411, 5414, 5419: oled_data = 16'b1111111100111101;
        5421, 5424, 5429, 5433, 5435, 5438, 5441, 5444, 5447, 5449: oled_data = 16'b1111111100111101;
        5453, 5454, 5456, 5458, 5459, 5461, 5462, 5464, 5466, 5469: oled_data = 16'b1111111100111101;
        5472, 5474, 5475, 5477, 5481, 5483, 5485, 5489, 5493, 5495: oled_data = 16'b1111111100111101;
        5499, 5501, 5503, 5506, 5508, 5510, 5512, 5513, 5515, 5516: oled_data = 16'b1111111100111101;
        5518, 5520, 5522, 5526, 5528, 5531, 5535, 5541, 5543, 5544: oled_data = 16'b1111111100111101;
        5546, 5547, 5549, 5551, 5553, 5555, 5560, 5563, 5568, 5578: oled_data = 16'b1111111100111101;
        5580, 5583, 5584, 5586, 5587, 5590, 5592, 5596, 5598, 5600: oled_data = 16'b1111111100111101;
        5603, 5607, 5609, 5615, 5617, 5619, 5620, 5622, 5629, 5631: oled_data = 16'b1111111100111101;
        5633, 5634, 5638, 5640, 5644, 5650, 5654, 5657, 5659, 5662: oled_data = 16'b1111111100111101;
        5663, 5666, 5669, 5673, 5675, 5677, 5681, 5684, 5689, 5691: oled_data = 16'b1111111100111101;
        5693, 5700, 5702, 5705, 5707, 5714, 5716, 5719, 5721, 5725: oled_data = 16'b1111111100111101;
        5728, 5730, 5732, 5737, 5739, 5741, 5744, 5747, 5751, 5753: oled_data = 16'b1111111100111101;
        5754, 5756, 5760, 5762, 5765, 5767, 5771, 5775, 5777, 5778: oled_data = 16'b1111111100111101;
        5781, 5783, 5786, 5790, 5792, 5793, 5796, 5799, 5801, 5802: oled_data = 16'b1111111100111101;
        5805, 5807, 5808, 5810, 5813, 5819, 5821, 5824, 5827, 5830: oled_data = 16'b1111111100111101;
        5833, 5835, 5836, 5838, 5839, 5841, 5844, 5847, 5849, 5854: oled_data = 16'b1111111100111101;
        5856, 5859, 5862, 5864, 5866, 5868, 5869, 5871, 5875, 5877: oled_data = 16'b1111111100111101;
        5878, 5880, 5883, 5899, 5901, 5902, 5907, 5911, 5918, 5920: oled_data = 16'b1111111100111101;
        5925, 5927, 5930, 5934, 5936, 5939, 5941, 5943, 5944, 5946: oled_data = 16'b1111111100111101;
        5948, 5951, 5961, 5966, 5968, 5972, 5974, 5975, 5977, 5980: oled_data = 16'b1111111100111101;
        5982, 5983, 5986, 5988, 5991, 5992, 5996, 5998, 6001, 6005: oled_data = 16'b1111111100111101;
        6008, 6010, 6011, 6014, 6018, 6022, 6025, 6027, 6029, 6031: oled_data = 16'b1111111100111101;
        6033, 6037, 6041, 6048, 6050, 6053, 6058, 6062, 6063, 6065: oled_data = 16'b1111111100111101;
        6066, 6072, 6074, 6080, 6082, 6083, 6085, 6089, 6091, 6095: oled_data = 16'b1111111100111101;
        6099, 6105, 6112, 6116, 6121, 6122, 6125, 6126, 6128, 6130: oled_data = 16'b1111111100111101;
        6132, 6134, 6135, 6137, 6140: oled_data = 16'b1111111100111101;
        1, 13, 16, 28, 31, 43, 46, 58, 61, 73: oled_data = 16'b1111011011111101;
        76, 88, 91, 107, 110, 122, 125, 137, 140, 152: oled_data = 16'b1111011011111101;
        
        155, 167, 170, 182, 185, 195, 198, 210, 213, 225: oled_data = 16'b1111011011111101;
        228, 240, 243, 255, 258, 270, 273, 285, 289, 292: oled_data = 16'b1111011011111101;
        300, 302, 310, 312, 320, 322, 330, 332, 340, 342: oled_data = 16'b1111011011111101;
        350, 352, 360, 362, 370, 372, 380, 391, 399, 411: oled_data = 16'b1111011011111101;
        439, 451, 459, 471, 488, 490, 493, 498, 520, 525: oled_data = 16'b1111011011111101;
        528, 530, 533, 538, 560, 565, 568, 570, 573, 579: oled_data = 16'b1111011011111101;
        594, 607, 612, 614, 617, 619, 637, 639, 642, 644: oled_data = 16'b1111011011111101;
        649, 662, 667, 669, 676, 691, 711, 716, 723, 736: oled_data = 16'b1111011011111101;
        743, 748, 769, 788, 790, 792, 797, 810, 815, 817: oled_data = 16'b1111011011111101;
        820, 822, 840, 842, 845, 847, 852, 868, 894, 901: oled_data = 16'b1111011011111101;
        904, 906, 924, 936, 946, 949, 954, 956, 963, 970: oled_data = 16'b1111011011111101;
        975, 989, 998, 1005, 1008, 1010, 1028, 1030, 1033, 1040: oled_data = 16'b1111011011111101;
        1053, 1057, 1072, 1076, 1084, 1087, 1090, 1114, 1119, 1122: oled_data = 16'b1111011011111101;
        1127, 1132, 1151, 1161, 1163, 1172, 1178, 1184, 1187, 1203: oled_data = 16'b1111011011111101;
        1213, 1216, 1221, 1223, 1241, 1257, 1262, 1276, 1281, 1284: oled_data = 16'b1111011011111101;
        1293, 1295, 1297, 1300, 1307, 1320, 1325, 1327, 1332, 1347: oled_data = 16'b1111011011111101;
        1351, 1356, 1424, 1431, 1444, 1449, 1520, 1530, 1537, 1547: oled_data = 16'b1111011011111101;
        1622, 1629, 1636, 1639, 1641, 1644, 1719, 1725, 1731, 1733: oled_data = 16'b1111011011111101;
        1738, 1741, 1812, 1816, 1825, 1909, 1928, 1931, 2009, 2020: oled_data = 16'b1111011011111101;
        2029, 2098, 2100, 2103, 2115, 2120, 2125, 2128, 2196, 2198: oled_data = 16'b1111011011111101;
        2202, 2220, 2299, 2302, 2305, 2311, 2319, 2321, 2336, 2347: oled_data = 16'b1111011011111101;
        2359, 2367, 2377, 2390, 2404, 2410, 2413, 2416, 2418, 2420: oled_data = 16'b1111011011111101;
        2422, 2427, 2444, 2456, 2467, 2474, 2487, 2492, 2499, 2510: oled_data = 16'b1111011011111101;
        2513, 2522, 2533, 2538, 2545, 2547, 2549, 2561, 2564, 2566: oled_data = 16'b1111011011111101;
        2578, 2586, 2589, 2593, 2596, 2598, 2610, 2622, 2630, 2632: oled_data = 16'b1111011011111101;
        2640, 2642, 2645, 2649, 2651, 2653, 2658, 2669, 2671, 2684: oled_data = 16'b1111011011111101;
        2697, 2699, 2701, 2704, 2707, 2710, 2731, 2742, 2759, 2761: oled_data = 16'b1111011011111101;
        2768, 2770, 2776, 2779, 2798, 2825, 2828, 2845, 2873, 2878: oled_data = 16'b1111011011111101;
        2881, 2883, 2885, 2892, 2912, 2920, 2922, 2925, 2957, 2966: oled_data = 16'b1111011011111101;
        2968, 2970, 2977, 2980, 2986, 3019, 3054, 3091, 3116, 3136: oled_data = 16'b1111011011111101;
        3148, 3160, 3162, 3164, 3198, 3211, 3233, 3255, 3258, 3261: oled_data = 16'b1111011011111101;
        3265, 3327, 3334, 3352, 3364, 3366, 3369, 3403, 3424, 3435: oled_data = 16'b1111011011111101;
        3466, 3521, 3535, 3541, 3567, 3569, 3585, 3587, 3599, 3621: oled_data = 16'b1111011011111101;
        3630, 3632, 3661, 3666, 3668, 3672, 3675, 3688, 3690, 3699: oled_data = 16'b1111011011111101;
        3718, 3720, 3731, 3734, 3737, 3745, 3759, 3769, 3772, 3776: oled_data = 16'b1111011011111101;
        3785, 3791, 3794, 3798, 3800, 3802, 3804, 3822, 3825, 3828: oled_data = 16'b1111011011111101;
        3834, 3857, 3862, 3869, 3873, 3879, 3882, 3888, 3897, 3901: oled_data = 16'b1111011011111101;
        3904, 3911, 3914, 3919, 3922, 3931, 3933, 3949, 3951, 3956: oled_data = 16'b1111011011111101;
        3961, 3966, 3968, 3970, 3974, 3976, 3979, 3983, 3985, 3988: oled_data = 16'b1111011011111101;
        3998, 4001, 4006, 4008, 4011, 4016, 4018, 4033, 4038, 4046: oled_data = 16'b1111011011111101;
        4048, 4050, 4055, 4073, 4078, 4089, 4091, 4124, 4137, 4139: oled_data = 16'b1111011011111101;
        4161, 4166, 4178, 4188, 4204, 4214, 4236, 4258, 4263, 4291: oled_data = 16'b1111011011111101;
        
        4309, 4317, 4327, 4329, 4360, 4396, 4410, 4414, 4421, 4428: oled_data = 16'b1111011011111101;
        4467, 4502, 4504, 4507, 4509, 4513, 4525, 4583, 4594, 4596: oled_data = 16'b1111011011111101;
        4601, 4606, 4638, 4645, 4647, 4683, 4693, 4695, 4697, 4703: oled_data = 16'b1111011011111101;
        4724, 4747, 4755, 4796, 4798, 4801, 4803, 4813, 4818, 4875: oled_data = 16'b1111011011111101;
        4881, 4883, 4885, 4890, 4893, 4900, 4903, 4910, 4915, 4927: oled_data = 16'b1111011011111101;
        4931, 4938, 4987, 4990, 4997, 5003, 5010, 5012, 5016, 5024: oled_data = 16'b1111011011111101;
        5032, 5051, 5089, 5104, 5107, 5109, 5123, 5126, 5129, 5131: oled_data = 16'b1111011011111101;
        5137, 5143, 5153, 5155, 5157, 5160, 5163, 5169, 5178, 5180: oled_data = 16'b1111011011111101;
        5182, 5185, 5190, 5214, 5234, 5237, 5240, 5257, 5262, 5266: oled_data = 16'b1111011011111101;
        5271, 5273, 5287, 5290, 5311, 5313, 5331, 5334, 5337, 5340: oled_data = 16'b1111011011111101;
        5345, 5351, 5356, 5358, 5366, 5379, 5387, 5403, 5410, 5420: oled_data = 16'b1111011011111101;
        5428, 5434, 5455, 5460, 5463, 5465, 5473, 5476, 5482, 5486: oled_data = 16'b1111011011111101;
        5488, 5500, 5502, 5509, 5514, 5519, 5527, 5545, 5548, 5550: oled_data = 16'b1111011011111101;
        5554, 5585, 5593, 5597, 5604, 5606, 5618, 5621, 5630, 5632: oled_data = 16'b1111011011111101;
        5637, 5639, 5649, 5658, 5676, 5682, 5690, 5706, 5715, 5729: oled_data = 16'b1111011011111101;
        5731, 5738, 5740, 5743, 5752, 5755, 5761, 5766, 5776, 5782: oled_data = 16'b1111011011111101;
        5791, 5800, 5803, 5806, 5809, 5820, 5837, 5840, 5848, 5850: oled_data = 16'b1111011011111101;
        5867, 5876, 5884, 5900, 5903, 5926, 5931, 5933, 5935, 5940: oled_data = 16'b1111011011111101;
        5945, 5967, 5973, 5976, 5984, 5987, 5993, 5997, 6009, 6030: oled_data = 16'b1111011011111101;
        6064, 6073, 6081, 6084, 6090, 6106, 6120, 6123, 6127, 6129: oled_data = 16'b1111011011111101;
        6133, 6136: oled_data = 16'b1111011011111101;
        3, 6, 8, 11, 18, 21, 23, 26, 33, 36: oled_data = 16'b1111111011111101;
        38, 41, 48, 51, 53, 56, 63, 66, 68, 71: oled_data = 16'b1111111011111101;
        78, 81, 83, 86, 93, 97, 100, 102, 105, 112: oled_data = 16'b1111111011111101;
        115, 117, 120, 127, 130, 132, 135, 142, 145, 147: oled_data = 16'b1111111011111101;
        150, 157, 160, 162, 165, 172, 175, 177, 180, 187: oled_data = 16'b1111111011111101;
        190, 193, 200, 203, 205, 208, 215, 218, 220, 223: oled_data = 16'b1111111011111101;
        230, 233, 235, 238, 245, 248, 250, 253, 260, 263: oled_data = 16'b1111111011111101;
        265, 268, 275, 278, 280, 283, 287, 295, 297, 305: oled_data = 16'b1111111011111101;
        307, 315, 317, 325, 327, 335, 337, 345, 347, 355: oled_data = 16'b1111111011111101;
        357, 365, 367, 375, 377, 385, 387, 389, 394, 396: oled_data = 16'b1111111011111101;
        406, 409, 414, 421, 424, 426, 429, 436, 441, 444: oled_data = 16'b1111111011111101;
        454, 456, 466, 469, 474, 478, 481, 484, 486, 495: oled_data = 16'b1111111011111101;
        500, 503, 505, 508, 510, 513, 515, 518, 523, 535: oled_data = 16'b1111111011111101;
        540, 543, 545, 548, 550, 553, 555, 558, 563, 575: oled_data = 16'b1111111011111101;
        577, 583, 586, 588, 590, 592, 597, 599, 602, 604: oled_data = 16'b1111111011111101;
        609, 622, 624, 627, 629, 632, 634, 647, 652, 654: oled_data = 16'b1111111011111101;
        657, 659, 664, 673, 677, 680, 683, 687, 693, 696: oled_data = 16'b1111111011111101;
        698, 701, 703, 706, 708, 713, 718, 721, 726, 728: oled_data = 16'b1111111011111101;
        731, 733, 738, 741, 746, 751, 753, 756, 758, 761: oled_data = 16'b1111111011111101;
        763, 766, 776, 780, 782, 784, 786, 795, 800, 802: oled_data = 16'b1111111011111101;
        805, 807, 812, 825, 827, 830, 832, 835, 837, 850: oled_data = 16'b1111111011111101;
        855, 857, 860, 862, 865, 870, 873, 876, 879, 889: oled_data = 16'b1111111011111101;
        891, 909, 916, 919, 921, 931, 934, 939, 951, 959: oled_data = 16'b1111111011111101;
        961, 966, 968, 973, 978, 981, 984, 987, 991, 993: oled_data = 16'b1111111011111101;
        
        995, 1000, 1003, 1013, 1015, 1018, 1020, 1023, 1025, 1035: oled_data = 16'b1111111011111101;
        1038, 1043, 1045, 1048, 1050, 1060, 1063, 1066, 1068, 1070: oled_data = 16'b1111111011111101;
        1074, 1078, 1081, 1092, 1094, 1097, 1099, 1102, 1104, 1107: oled_data = 16'b1111111011111101;
        1109, 1112, 1117, 1124, 1129, 1134, 1137, 1139, 1142, 1144: oled_data = 16'b1111111011111101;
        1147, 1149, 1153, 1155, 1157, 1159, 1166, 1180, 1182, 1190: oled_data = 16'b1111111011111101;
        1192, 1194, 1196, 1198, 1201, 1206, 1208, 1211, 1218, 1226: oled_data = 16'b1111111011111101;
        1228, 1231, 1233, 1236, 1238, 1243, 1246, 1249, 1252, 1254: oled_data = 16'b1111111011111101;
        1260, 1279, 1287, 1290, 1302, 1305, 1310, 1312, 1315, 1317: oled_data = 16'b1111111011111101;
        1322, 1330, 1335, 1337, 1340, 1342, 1345, 1354, 1434, 1436: oled_data = 16'b1111111011111101;
        1439, 1441, 1445, 1447, 1452, 1522, 1524, 1526, 1528, 1533: oled_data = 16'b1111111011111101;
        1539, 1542, 1545, 1619, 1625, 1627, 1631, 1633, 1714, 1716: oled_data = 16'b1111111011111101;
        1722, 1729, 1735, 1814, 1819, 1823, 1831, 1833, 1835, 1837: oled_data = 16'b1111111011111101;
        1906, 1912, 1914, 1916, 1918, 1921, 1923, 1925, 1934, 2003: oled_data = 16'b1111111011111101;
        2005, 2007, 2012, 2015, 2017, 2022, 2025, 2027, 2106, 2109: oled_data = 16'b1111111011111101;
        2113, 2118, 2122, 2127, 2193, 2200, 2204, 2206, 2209, 2212: oled_data = 16'b1111111011111101;
        2215, 2218, 2225, 2287, 2290, 2293, 2296, 2307, 2309, 2313: oled_data = 16'b1111111011111101;
        2316, 2318, 2323, 2327, 2330, 2332, 2334, 2337, 2339, 2341: oled_data = 16'b1111111011111101;
        2343, 2345, 2349, 2351, 2353, 2355, 2357, 2361, 2363, 2365: oled_data = 16'b1111111011111101;
        2369, 2371, 2373, 2375, 2379, 2381, 2384, 2386, 2388, 2393: oled_data = 16'b1111111011111101;
        2395, 2397, 2399, 2401, 2407, 2424, 2430, 2434, 2436, 2439: oled_data = 16'b1111111011111101;
        2442, 2446, 2448, 2451, 2454, 2458, 2461, 2463, 2465, 2470: oled_data = 16'b1111111011111101;
        2472, 2476, 2478, 2480, 2482, 2485, 2489, 2497, 2504, 2506: oled_data = 16'b1111111011111101;
        2517, 2520, 2524, 2527, 2528, 2531, 2536, 2541, 2552, 2555: oled_data = 16'b1111111011111101;
        2558, 2569, 2572, 2575, 2580, 2583, 2590, 2600, 2603, 2606: oled_data = 16'b1111111011111101;
        2608, 2612, 2614, 2617, 2620, 2625, 2628, 2635, 2638, 2647: oled_data = 16'b1111111011111101;
        2655, 2660, 2663, 2666, 2676, 2680, 2682, 2687, 2689, 2691: oled_data = 16'b1111111011111101;
        2694, 2712, 2714, 2716, 2719, 2721, 2723, 2726, 2729, 2733: oled_data = 16'b1111111011111101;
        2735, 2738, 2740, 2745, 2748, 2751, 2753, 2755, 2757, 2763: oled_data = 16'b1111111011111101;
        2765, 2773, 2781, 2785, 2788, 2791, 2793, 2796, 2801, 2811: oled_data = 16'b1111111011111101;
        2834, 2839, 2860, 2862, 2865, 2867, 2870, 2875, 2887, 2890: oled_data = 16'b1111111011111101;
        2895, 2906, 2914, 2943, 2951, 2959, 2962, 2964, 2972, 2974: oled_data = 16'b1111111011111101;
        2984, 2989, 2993, 2994, 3021, 3023, 3051, 3056, 3059, 3062: oled_data = 16'b1111111011111101;
        3065, 3069, 3071, 3073, 3079, 3082, 3084, 3086, 3088, 3110: oled_data = 16'b1111111011111101;
        3131, 3143, 3151, 3153, 3156, 3158, 3169, 3172, 3173, 3176: oled_data = 16'b1111111011111101;
        3179, 3183, 3185, 3187, 3192, 3214, 3231, 3237, 3243, 3245: oled_data = 16'b1111111011111101;
        3248, 3250, 3252, 3262, 3267, 3270, 3272, 3274, 3276, 3278: oled_data = 16'b1111111011111101;
        3282, 3289, 3294, 3307, 3309, 3319, 3340, 3342, 3345, 3348: oled_data = 16'b1111111011111101;
        3350, 3359, 3361, 3372, 3375, 3376, 3379, 3406, 3429, 3431: oled_data = 16'b1111111011111101;
        3440, 3442, 3444, 3447, 3451, 3453, 3455, 3457, 3459, 3462: oled_data = 16'b1111111011111101;
        3469, 3473, 3481, 3500, 3502, 3526, 3531, 3533, 3544, 3547: oled_data = 16'b1111111011111101;
        3549, 3553, 3556, 3559, 3562, 3564, 3571, 3578, 3594, 3596: oled_data = 16'b1111111011111101;
        
        3608, 3615, 3617, 3627, 3635, 3637, 3639, 3641, 3644, 3646: oled_data = 16'b1111111011111101;
        3649, 3651, 3653, 3655, 3657, 3659, 3664, 3682, 3684, 3693: oled_data = 16'b1111111011111101;
        3696, 3705, 3711, 3714, 3724, 3727, 3729, 3739, 3748, 3750: oled_data = 16'b1111111011111101;
        3753, 3756, 3763, 3767, 3779, 3782, 3787, 3789, 3806, 3808: oled_data = 16'b1111111011111101;
        3811, 3813, 3816, 3818, 3820, 3830, 3832, 3836, 3839, 3841: oled_data = 16'b1111111011111101;
        3843, 3847, 3850, 3853, 3856, 3860, 3865, 3867, 3871, 3876: oled_data = 16'b1111111011111101;
        3885, 3890, 3892, 3894, 3906, 3909, 3917, 3924, 3927, 3937: oled_data = 16'b1111111011111101;
        3940, 3941, 3945, 3947, 3959, 3972, 3981, 3991, 3994, 3996: oled_data = 16'b1111111011111101;
        4003, 4014, 4021, 4024, 4029, 4031, 4035, 4041, 4044, 4053: oled_data = 16'b1111111011111101;
        4061, 4068, 4071, 4075, 4081, 4083, 4085, 4094, 4096, 4101: oled_data = 16'b1111111011111101;
        4104, 4106, 4108, 4111, 4114, 4116, 4118, 4120, 4122, 4129: oled_data = 16'b1111111011111101;
        4135, 4148, 4169, 4172, 4186, 4199, 4205, 4208, 4211, 4217: oled_data = 16'b1111111011111101;
        4220, 4223, 4225, 4227, 4229, 4231, 4256, 4265, 4275, 4299: oled_data = 16'b1111111011111101;
        4301, 4305, 4307, 4314, 4321, 4324, 4358, 4363, 4379, 4391: oled_data = 16'b1111111011111101;
        4397, 4402, 4405, 4408, 4412, 4417, 4424, 4426, 4455, 4457: oled_data = 16'b1111111011111101;
        4463, 4499, 4511, 4516, 4518, 4521, 4523, 4549, 4552, 4554: oled_data = 16'b1111111011111101;
        4571, 4598, 4603, 4609, 4611, 4614, 4616, 4620, 4650, 4659: oled_data = 16'b1111111011111101;
        4689, 4691, 4700, 4705, 4708, 4711, 4713, 4715, 4717, 4740: oled_data = 16'b1111111011111101;
        4745, 4763, 4775, 4785, 4788, 4791, 4794, 4805, 4807, 4837: oled_data = 16'b1111111011111101;
        4840, 4851, 4863, 4888, 4895, 4897, 4905, 4907, 4934, 4936: oled_data = 16'b1111111011111101;
        4943, 4955, 4959, 4963, 4973, 4977, 4981, 4983, 4985, 4993: oled_data = 16'b1111111011111101;
        4995, 5000, 5021, 5029, 5040, 5044, 5055, 5068, 5074, 5076: oled_data = 16'b1111111011111101;
        5079, 5083, 5085, 5092, 5094, 5097, 5099, 5102, 5111, 5113: oled_data = 16'b1111111011111101;
        5115, 5117, 5119, 5122, 5133, 5139, 5141, 5145, 5148, 5150: oled_data = 16'b1111111011111101;
        5159, 5165, 5167, 5171, 5173, 5176, 5192, 5194, 5196, 5198: oled_data = 16'b1111111011111101;
        5200, 5202, 5205, 5208, 5211, 5216, 5220, 5222, 5227, 5230: oled_data = 16'b1111111011111101;
        5232, 5242, 5244, 5246, 5248, 5251, 5253, 5259, 5276, 5279: oled_data = 16'b1111111011111101;
        5281, 5284, 5293, 5296, 5299, 5302, 5305, 5308, 5317, 5319: oled_data = 16'b1111111011111101;
        5321, 5324, 5326, 5329, 5343, 5348, 5350, 5353, 5360, 5362: oled_data = 16'b1111111011111101;
        5364, 5369, 5371, 5373, 5377, 5381, 5383, 5385, 5390, 5393: oled_data = 16'b1111111011111101;
        5395, 5397, 5399, 5401, 5405, 5408, 5412, 5416, 5418, 5423: oled_data = 16'b1111111011111101;
        5426, 5430, 5432, 5437, 5440, 5442, 5445, 5450, 5452, 5457: oled_data = 16'b1111111011111101;
        5468, 5470, 5479, 5484, 5490, 5492, 5496, 5498, 5505, 5511: oled_data = 16'b1111111011111101;
        5524, 5530, 5534, 5537, 5539, 5557, 5559, 5562, 5567, 5569: oled_data = 16'b1111111011111101;
        5573, 5576, 5582, 5589, 5602, 5611, 5613, 5616, 5623, 5625: oled_data = 16'b1111111011111101;
        5627, 5635, 5642, 5645, 5647, 5653, 5660, 5665, 5668, 5670: oled_data = 16'b1111111011111101;
        5672, 5674, 5679, 5683, 5686, 5688, 5692, 5695, 5697, 5701: oled_data = 16'b1111111011111101;
        5704, 5708, 5710, 5712, 5717, 5720, 5724, 5726, 5734, 5736: oled_data = 16'b1111111011111101;
        5745, 5748, 5750, 5757, 5759, 5763, 5769, 5772, 5774, 5780: oled_data = 16'b1111111011111101;
        5784, 5787, 5789, 5794, 5798, 5811, 5816, 5818, 5823, 5825: oled_data = 16'b1111111011111101;
        5828, 5831, 5834, 5842, 5845, 5853, 5857, 5860, 5863, 5872: oled_data = 16'b1111111011111101;
        
        5881, 5887, 5889, 5891, 5893, 5895, 5897, 5905, 5908, 5910: oled_data = 16'b1111111011111101;
        5913, 5915, 5917, 5922, 5924, 5928, 5938, 5947, 5950, 5953: oled_data = 16'b1111111011111101;
        5955, 5957, 5962, 5964, 5969, 5971, 5978, 5981, 5989, 5995: oled_data = 16'b1111111011111101;
        5999, 6002, 6007, 6012, 6015, 6017, 6021, 6024, 6028, 6032: oled_data = 16'b1111111011111101;
        6035, 6038, 6040, 6043, 6045, 6047, 6049, 6052, 6054, 6056: oled_data = 16'b1111111011111101;
        6059, 6061, 6068, 6070, 6075, 6077, 6079, 6086, 6088, 6093: oled_data = 16'b1111111011111101;
        6096, 6098, 6101, 6103, 6109, 6111, 6114, 6118, 6138, 6141: oled_data = 16'b1111111011111101;
        4, 7, 10, 19, 22, 25, 34, 37, 40, 49: oled_data = 16'b1111011100111101;
        52, 55, 64, 67, 70, 79, 82, 85, 94, 98: oled_data = 16'b1111011100111101;
        101, 104, 113, 116, 119, 128, 131, 134, 143, 146: oled_data = 16'b1111011100111101;
        149, 158, 161, 164, 173, 176, 179, 188, 191, 192: oled_data = 16'b1111011100111101;
        201, 204, 207, 216, 219, 222, 231, 234, 237, 246: oled_data = 16'b1111011100111101;
        249, 252, 261, 264, 267, 276, 279, 282, 294, 296: oled_data = 16'b1111011100111101;
        298, 304, 306, 308, 314, 316, 318, 324, 326, 328: oled_data = 16'b1111011100111101;
        334, 336, 338, 344, 346, 348, 354, 356, 358, 364: oled_data = 16'b1111011100111101;
        366, 368, 374, 376, 378, 382, 386, 403, 415, 423: oled_data = 16'b1111011100111101;
        427, 435, 447, 463, 475, 479, 480, 482, 485, 496: oled_data = 16'b1111011100111101;
        501, 504, 506, 509, 512, 514, 517, 522, 536, 541: oled_data = 16'b1111011100111101;
        544, 546, 549, 552, 554, 557, 562, 582, 585, 587: oled_data = 16'b1111011100111101;
        589, 591, 596, 598, 601, 603, 605, 610, 621, 623: oled_data = 16'b1111011100111101;
        626, 628, 630, 633, 635, 646, 651, 653, 655, 658: oled_data = 16'b1111011100111101;
        660, 665, 671, 672, 674, 679, 684, 688, 695, 700: oled_data = 16'b1111011100111101;
        704, 707, 720, 727, 732, 739, 752, 755, 759, 764: oled_data = 16'b1111011100111101;
        773, 775, 777, 781, 783, 785, 794, 799, 801, 804: oled_data = 16'b1111011100111101;
        806, 808, 813, 824, 826, 829, 831, 833, 836, 838: oled_data = 16'b1111011100111101;
        849, 854, 856, 858, 863, 866, 872, 875, 882, 885: oled_data = 16'b1111011100111101;
        888, 892, 898, 910, 922, 930, 933, 940, 942, 952: oled_data = 16'b1111011100111101;
        958, 960, 965, 967, 972, 977, 979, 982, 985, 992: oled_data = 16'b1111011100111101;
        994, 996, 1001, 1012, 1014, 1017, 1021, 1024, 1026, 1037: oled_data = 16'b1111011100111101;
        1042, 1044, 1046, 1049, 1061, 1064, 1069, 1079, 1082, 1095: oled_data = 16'b1111011100111101;
        1098, 1100, 1103, 1106, 1111, 1116, 1130, 1135, 1138, 1143: oled_data = 16'b1111011100111101;
        1146, 1148, 1154, 1158, 1165, 1181, 1189, 1191, 1193, 1197: oled_data = 16'b1111011100111101;
        1200, 1205, 1207, 1209, 1219, 1225, 1229, 1232, 1235, 1237: oled_data = 16'b1111011100111101;
        1239, 1248, 1250, 1255, 1259, 1278, 1288, 1291, 1304, 1309: oled_data = 16'b1111011100111101;
        1311, 1313, 1316, 1323, 1329, 1336, 1339, 1341, 1343, 1349: oled_data = 16'b1111011100111101;
        1433, 1435, 1438, 1440, 1442, 1446, 1450, 1523, 1525, 1532: oled_data = 16'b1111011100111101;
        1535, 1541, 1618, 1624, 1634, 1715, 1717, 1721, 1723, 1727: oled_data = 16'b1111011100111101;
        1728, 1818, 1822, 1830, 1832, 1834, 1838, 1846, 1907, 1917: oled_data = 16'b1111011100111101;
        1922, 1924, 1926, 2006, 2011, 2014, 2016, 2018, 2023, 2031: oled_data = 16'b1111011100111101;
        2105, 2108, 2111, 2117, 2123, 2191, 2194, 2205, 2208, 2210: oled_data = 16'b1111011100111101;
        2214, 2217, 2222, 2288, 2292, 2295, 2297, 2308, 2314, 2328: oled_data = 16'b1111011100111101;
        2333, 2340, 2344, 2350, 2352, 2354, 2356, 2362, 2364, 2370: oled_data = 16'b1111011100111101;
        2372, 2374, 2380, 2383, 2385, 2396, 2398, 2402, 2406, 2408: oled_data = 16'b1111011100111101;
        2412, 2425, 2429, 2431, 2433, 2435, 2438, 2441, 2447, 2453: oled_data = 16'b1111011100111101;
        
        2459, 2462, 2464, 2471, 2477, 2481, 2484, 2490, 2495, 2496: oled_data = 16'b1111011100111101;
        2503, 2507, 2516, 2519, 2525, 2530, 2535, 2540, 2542, 2551: oled_data = 16'b1111011100111101;
        2553, 2556, 2559, 2568, 2571, 2574, 2576, 2581, 2584, 2601: oled_data = 16'b1111011100111101;
        2604, 2607, 2613, 2616, 2619, 2624, 2627, 2634, 2637, 2661: oled_data = 16'b1111011100111101;
        2665, 2667, 2675, 2681, 2686, 2690, 2693, 2695, 2713, 2715: oled_data = 16'b1111011100111101;
        2717, 2720, 2722, 2724, 2728, 2734, 2737, 2739, 2744, 2750: oled_data = 16'b1111011100111101;
        2752, 2754, 2756, 2764, 2772, 2774, 2783, 2784, 2787, 2792: oled_data = 16'b1111011100111101;
        2800, 2809, 2818, 2847, 2855, 2861, 2863, 2866, 2869, 2876: oled_data = 16'b1111011100111101;
        2886, 2889, 2891, 2894, 2897, 2907, 2915, 2936, 2955, 2960: oled_data = 16'b1111011100111101;
        2963, 2973, 2983, 3022, 3047, 3057, 3067, 3070, 3074, 3077: oled_data = 16'b1111011100111101;
        3080, 3083, 3087, 3089, 3127, 3142, 3150, 3152, 3157, 3167: oled_data = 16'b1111011100111101;
        3168, 3171, 3174, 3177, 3180, 3184, 3193, 3197, 3206, 3215: oled_data = 16'b1111011100111101;
        3244, 3247, 3251, 3253, 3268, 3271, 3273, 3275, 3277, 3279: oled_data = 16'b1111011100111101;
        3281, 3283, 3288, 3293, 3308, 3310, 3341, 3344, 3346, 3349: oled_data = 16'b1111011100111101;
        3358, 3362, 3373, 3377, 3389, 3390, 3407, 3415, 3419, 3430: oled_data = 16'b1111011100111101;
        3441, 3443, 3446, 3452, 3454, 3456, 3458, 3461, 3463, 3468: oled_data = 16'b1111011100111101;
        3470, 3475, 3480, 3498, 3501, 3527, 3532, 3539, 3546, 3548: oled_data = 16'b1111011100111101;
        3551, 3555, 3560, 3563, 3577, 3593, 3595, 3597, 3607, 3616: oled_data = 16'b1111011100111101;
        3628, 3634, 3640, 3642, 3645, 3648, 3650, 3652, 3654, 3656: oled_data = 16'b1111011100111101;
        3658, 3681, 3683, 3694, 3704, 3710, 3713, 3725, 3728, 3733: oled_data = 16'b1111011100111101;
        3740, 3749, 3752, 3755, 3757, 3760, 3762, 3765, 3774, 3780: oled_data = 16'b1111011100111101;
        3788, 3807, 3810, 3812, 3814, 3817, 3819, 3831, 3838, 3842: oled_data = 16'b1111011100111101;
        3844, 3846, 3849, 3852, 3859, 3864, 3866, 3875, 3877, 3884: oled_data = 16'b1111011100111101;
        3886, 3891, 3893, 3907, 3916, 3925, 3928, 3936, 3939, 3946: oled_data = 16'b1111011100111101;
        3958, 3963, 3990, 3992, 3995, 4004, 4013, 4020, 4022, 4025: oled_data = 16'b1111011100111101;
        4027, 4030, 4036, 4040, 4043, 4052, 4060, 4063, 4067, 4069: oled_data = 16'b1111011100111101;
        4076, 4082, 4086, 4093, 4097, 4102, 4105, 4110, 4112, 4115: oled_data = 16'b1111011100111101;
        4119, 4121, 4127, 4130, 4133, 4154, 4168, 4170, 4180, 4185: oled_data = 16'b1111011100111101;
        4194, 4212, 4218, 4221, 4224, 4226, 4228, 4230, 4232, 4244: oled_data = 16'b1111011100111101;
        4276, 4282, 4300, 4306, 4313, 4315, 4319, 4323, 4331, 4362: oled_data = 16'b1111011100111101;
        4403, 4407, 4416, 4418, 4425, 4430, 4435, 4436, 4454, 4456: oled_data = 16'b1111011100111101;
        4459, 4483, 4497, 4500, 4515, 4517, 4519, 4522, 4526, 4530: oled_data = 16'b1111011100111101;
        4531, 4540, 4541, 4548, 4553, 4604, 4612, 4615, 4617, 4619: oled_data = 16'b1111011100111101;
        4622, 4627, 4636, 4643, 4649, 4651, 4690, 4699, 4704, 4706: oled_data = 16'b1111011100111101;
        4709, 4712, 4716, 4718, 4722, 4732, 4734, 4735, 4739, 4741: oled_data = 16'b1111011100111101;
        4744, 4787, 4790, 4793, 4806, 4809, 4811, 4819, 4820, 4824: oled_data = 16'b1111011100111101;
        4828, 4829, 4830, 4831, 4835, 4836, 4838, 4841, 4847, 4887: oled_data = 16'b1111011100111101;
        4898, 4906, 4914, 4916, 4920, 4924, 4925, 4926, 4933, 4935: oled_data = 16'b1111011100111101;
        4947, 4978, 4982, 4984, 4992, 4999, 5001, 5007, 5020, 5022: oled_data = 16'b1111011100111101;
        5023, 5027, 5028, 5035, 5039, 5043, 5045, 5063, 5067, 5069: oled_data = 16'b1111011100111101;
        5075, 5077, 5081, 5084, 5087, 5091, 5093, 5096, 5100, 5112: oled_data = 16'b1111011100111101;
        
        5114, 5116, 5120, 5121, 5134, 5140, 5146, 5149, 5151, 5172: oled_data = 16'b1111011100111101;
        5193, 5197, 5199, 5201, 5204, 5206, 5209, 5212, 5218, 5221: oled_data = 16'b1111011100111101;
        5223, 5225, 5228, 5231, 5243, 5247, 5250, 5254, 5260, 5264: oled_data = 16'b1111011100111101;
        5277, 5282, 5285, 5294, 5298, 5301, 5303, 5306, 5309, 5316: oled_data = 16'b1111011100111101;
        5320, 5323, 5325, 5328, 5342, 5347, 5349, 5361, 5363, 5370: oled_data = 16'b1111011100111101;
        5372, 5374, 5376, 5384, 5389, 5392, 5394, 5396, 5400, 5407: oled_data = 16'b1111011100111101;
        5413, 5415, 5417, 5422, 5425, 5436, 5439, 5443, 5446, 5451: oled_data = 16'b1111011100111101;
        5467, 5471, 5478, 5480, 5497, 5504, 5507, 5523, 5525, 5529: oled_data = 16'b1111011100111101;
        5533, 5538, 5540, 5552, 5556, 5558, 5561, 5564, 5566, 5570: oled_data = 16'b1111011100111101;
        5572, 5574, 5577, 5581, 5588, 5591, 5595, 5601, 5610, 5612: oled_data = 16'b1111011100111101;
        5614, 5624, 5626, 5628, 5641, 5643, 5646, 5652, 5655, 5661: oled_data = 16'b1111011100111101;
        5664, 5667, 5671, 5678, 5680, 5685, 5687, 5694, 5696, 5698: oled_data = 16'b1111011100111101;
        5703, 5709, 5711, 5713, 5718, 5723, 5727, 5733, 5735, 5746: oled_data = 16'b1111011100111101;
        5749, 5758, 5764, 5768, 5770, 5773, 5779, 5785, 5788, 5795: oled_data = 16'b1111011100111101;
        5797, 5812, 5815, 5817, 5822, 5826, 5829, 5832, 5843, 5846: oled_data = 16'b1111011100111101;
        5852, 5855, 5858, 5861, 5873, 5882, 5886, 5888, 5890, 5892: oled_data = 16'b1111011100111101;
        5894, 5896, 5898, 5906, 5909, 5912, 5914, 5916, 5921, 5923: oled_data = 16'b1111011100111101;
        5929, 5937, 5949, 5952, 5954, 5958, 5960, 5963, 5965, 5970: oled_data = 16'b1111011100111101;
        5990, 6000, 6003, 6006, 6016, 6020, 6023, 6034, 6036, 6039: oled_data = 16'b1111011100111101;
        6042, 6044, 6046, 6051, 6055, 6057, 6060, 6067, 6069, 6071: oled_data = 16'b1111011100111101;
        6076, 6078, 6092, 6094, 6097, 6100, 6102, 6104, 6108, 6110: oled_data = 16'b1111011100111101;
        6113, 6115, 6117, 6124, 6139, 6143: oled_data = 16'b1111011100111101;
        388, 395, 407, 443, 455, 467, 861, 878, 890, 908: oled_data = 16'b1111011100111100;
        917, 920, 938, 1156, 1167, 1173, 1245, 1357, 1544, 1836: oled_data = 16'b1111011100111100;
        1911, 1915, 2026, 2387, 2392, 3060, 3063, 3085, 3154, 3472: oled_data = 16'b1111011100111100;
        3543, 4095, 4209, 5175, 5195, 5354, 5431, 5491, 5536, 5956: oled_data = 16'b1111011100111100;
        5979, 6013, 6087: oled_data = 16'b1111011100111100;
        392, 398, 410, 413, 422, 425, 428, 437, 440, 452: oled_data = 16'b1111111100111100;
        458, 470, 473, 893, 902, 905, 923, 932, 935, 947: oled_data = 16'b1111111100111100;
        950, 953, 1160, 1164, 1338, 1423, 1432, 1443, 1734, 2101: oled_data = 16'b1111111100111100;
        2211, 2216, 2298, 2414, 2417, 2494, 2595, 2602, 2741, 2767: oled_data = 16'b1111111100111100;
        2780, 2826, 2835, 2874, 2888, 3053, 3370, 3404, 3460, 3747: oled_data = 16'b1111111100111100;
        3786, 3790, 3823, 3829, 3851, 3880, 3923, 3971, 3993, 4047: oled_data = 16'b1111111100111100;
        4103, 4107, 4179, 4328, 4361, 4411, 4501, 4701, 4710, 4792: oled_data = 16'b1111111100111100;
        4795, 4804, 4884, 5191, 5261, 5265, 5275, 5427, 5487, 5575: oled_data = 16'b1111111100111100;
        5594, 5605, 5636, 5648, 5722, 5742, 5804, 5851, 5885, 5904: oled_data = 16'b1111111100111100;
        5932, 5985, 5994, 6107, 6119, 6142: oled_data = 16'b1111111100111100;
        401, 404, 416, 434, 446, 449, 461, 464, 476, 771: oled_data = 16'b1111111011111100;
        774, 881, 884, 887, 896, 899, 911, 929, 941, 944: oled_data = 16'b1111111011111100;
        1821, 1828, 2501, 2508, 2673, 2817, 2982, 3075, 3464, 3538: oled_data = 16'b1111111011111100;
        3566, 3954, 3964, 4026, 4058, 4065, 4087, 4126, 4132, 4193: oled_data = 16'b1111111011111100;
        4234, 4419, 4743, 4810, 4932, 4967, 5034, 5224, 5315, 5517: oled_data = 16'b1111111011111100;
        5532, 5542, 5565, 5571, 5599, 5651, 5656, 5699, 5814, 5874: oled_data = 16'b1111111011111100;
        
        5959, 6004, 6019, 6131: oled_data = 16'b1111111011111100;
        419, 431, 778, 914, 926, 1168, 1169, 1170, 1171, 1174: oled_data = 16'b1111011011111100;
        1175, 1176, 1177, 1426, 1429, 1453, 1549, 1645, 2678, 2831: oled_data = 16'b1111011011111100;
        2991, 3118, 3355, 3438, 3449, 3742, 3943, 4099, 4202, 4267: oled_data = 16'b1111011011111100;
        4311, 5005, 5187, 5269, 5448, 5494, 5521, 5579, 5608, 5865: oled_data = 16'b1111011011111100;
        5870, 5879, 5919, 5942, 6026: oled_data = 16'b1111011011111100;
        1263, 1839: oled_data = 16'b1001110001010011;
        1264, 1265, 1267, 1270, 1271, 1273, 1454, 1467, 1569, 1615: oled_data = 16'b0011100111001010;
        1646, 1762, 1808, 1840, 2049, 2131, 2134, 2136, 2138, 2140: oled_data = 16'b0011100111001010;
        2141, 2145, 2147, 2148, 2149, 2150, 2151, 2152, 2154, 2155: oled_data = 16'b0011100111001010;
        2156, 2157, 2158, 2159, 2160, 2161, 2162, 2163, 2164, 2165: oled_data = 16'b0011100111001010;
        2166, 2167, 2169, 2170, 2171, 2172, 2173, 2174, 2175, 2176: oled_data = 16'b0011100111001010;
        2177, 2179, 2180, 2181, 2182, 2183, 2184, 2186, 2187, 2188: oled_data = 16'b0011100111001010;
        2189: oled_data = 16'b0011100111001010;
        1266: oled_data = 16'b0011001000001010;
        1268: oled_data = 16'b1101110111111000;
        1269: oled_data = 16'b1011010011110101;
        1272, 2139, 2142: oled_data = 16'b0011000111001010;
        1274: oled_data = 16'b1011110100110101;
        1358, 1371, 1372, 1374, 1377, 1380, 1384, 1387, 1389, 1392: oled_data = 16'b1000001111010001;
        1393, 1395, 1396, 1398, 1401, 1404, 1405, 1407, 1408, 1411: oled_data = 16'b1000001111010001;
        1414, 1416, 1417, 1419, 1420: oled_data = 16'b1000001111010001;
        1359: oled_data = 16'b1000101100001110;
        1360, 2133: oled_data = 16'b1010001010001010;
        1361: oled_data = 16'b1010101100001100;
        1362, 1363, 1366, 1367, 1368, 1369: oled_data = 16'b1011001100001100;
        1364: oled_data = 16'b0111101110001111;
        1365: oled_data = 16'b1000101101001111;
        1370: oled_data = 16'b1000001101001111;
        1373, 1376, 1379, 1382, 1385, 1388, 1391, 1400, 1403, 1409: oled_data = 16'b1000001111010000;
        1412, 1421: oled_data = 16'b1000001111010000;
        1375, 1378, 1383, 1386, 1390, 1399, 1402, 1410, 1413: oled_data = 16'b0111101111010001;
        1381: oled_data = 16'b0111101110010001;
        1394, 1397, 1406, 1415, 1418: oled_data = 16'b0111101111010000;
        1422: oled_data = 16'b1011110101110111;
        1455, 1551, 1647: oled_data = 16'b1000001001001010;
        1456, 1648, 1939: oled_data = 16'b1101101011001010;
        1457, 1458, 1553, 1651, 1653: oled_data = 16'b1111101110001101;
        1459, 1555, 1652, 1749: oled_data = 16'b1111101111001110;
        1460: oled_data = 16'b0110001000001010;
        1461: oled_data = 16'b1000001010001011;
        1462, 1465, 1554, 1556, 1558, 1654, 1657, 1748: oled_data = 16'b1111101111001101;
        1463: oled_data = 16'b1111101111001111;
        1464: oled_data = 16'b1111110000001111;
        1466, 1755, 2228: oled_data = 16'b0110101001001010;
        1468, 1470, 1476, 1478, 1480, 1482, 1485, 1487, 1489, 1491: oled_data = 16'b0100101000001010;
        1494, 1496, 1498, 1500, 1503, 1505, 1507, 1509, 1512, 1514: oled_data = 16'b0100101000001010;
        1516: oled_data = 16'b0100101000001010;
        1469, 1471, 1659, 2039, 2095: oled_data = 16'b0101001000001010;
        1472: oled_data = 16'b0100000111001010;
        1473, 1904, 2135, 2143, 2146, 2153, 2168, 2178, 2185: oled_data = 16'b0011100111001001;
        1474, 1475, 1479, 1481, 1483, 1484, 1486, 1488, 1490, 1492: oled_data = 16'b0100101000001011;
        1493, 1495, 1497, 1499, 1501, 1502, 1504, 1506, 1508, 1510: oled_data = 16'b0100101000001011;
        1511, 1513, 1515, 1517: oled_data = 16'b0100101000001011;
        1477: oled_data = 16'b0100101001001011;
        1518, 2051, 2052, 2053, 2055, 2056, 2058, 2059, 2060, 2061: oled_data = 16'b1000101111010001;
        2063, 2064, 2065, 2066, 2067, 2068, 2070, 2071, 2073, 2074: oled_data = 16'b1000101111010001;
        2075, 2076, 2077, 2078, 2080, 2081, 2083, 2084, 2085, 2087: oled_data = 16'b1000101111010001;
        
        2088, 2090, 2091, 2093: oled_data = 16'b1000101111010001;
        1519: oled_data = 16'b1110011000111001;
        1550, 1849, 2137, 2144: oled_data = 16'b0011101000001010;
        1552, 1745, 1842: oled_data = 16'b1101101011001011;
        1557, 1561: oled_data = 16'b1111101110001110;
        1559: oled_data = 16'b1111011000111001;
        1560: oled_data = 16'b1111111001111001;
        1562: oled_data = 16'b0110001001001010;
        1563, 2040: oled_data = 16'b0101101000001010;
        1564, 1566, 1757, 1759, 1760, 1851, 1947, 1948, 1949, 1951: oled_data = 16'b1110101011001000;
        1565, 1567, 1756, 1853, 1855: oled_data = 16'b1110101011000111;
        1568: oled_data = 16'b0111101001001001;
        1570, 1573, 1579, 1581, 1586, 1588, 1591, 1596, 1598, 1602: oled_data = 16'b1010010010110100;
        1606, 1608, 1613, 1670, 1674, 1678, 1680, 1685, 1688, 1695: oled_data = 16'b1010010010110100;
        1697, 1700, 1703, 1706, 1764, 1767, 1772, 1779, 1782, 1785: oled_data = 16'b1010010010110100;
        1787, 1789, 1792, 1795, 1800, 1803, 1861, 1874, 1876, 1884: oled_data = 16'b1010010010110100;
        1889, 1894, 1900, 1902, 1958, 1963, 1966, 1968, 1976, 1983: oled_data = 16'b1010010010110100;
        1986, 1988, 1991, 1994, 1997, 2130: oled_data = 16'b1010010010110100;
        1571, 1572, 1574, 1575, 1576, 1577, 1578, 1580, 1582, 1583: oled_data = 16'b1010010010110101;
        1584, 1585, 1587, 1589, 1590, 1592, 1593, 1594, 1595, 1597: oled_data = 16'b1010010010110101;
        1599, 1600, 1601, 1603, 1604, 1605, 1607, 1609, 1610, 1611: oled_data = 16'b1010010010110101;
        1612, 1668, 1671, 1673, 1675, 1676, 1679, 1681, 1682, 1684: oled_data = 16'b1010010010110101;
        1686, 1689, 1691, 1692, 1694, 1698, 1701, 1704, 1707, 1709: oled_data = 16'b1010010010110101;
        1765, 1766, 1768, 1769, 1771, 1773, 1774, 1776, 1778, 1780: oled_data = 16'b1010010010110101;
        1783, 1784, 1786, 1790, 1791, 1793, 1794, 1796, 1798, 1799: oled_data = 16'b1010010010110101;
        1801, 1802, 1804, 1805, 1807, 1860, 1863, 1865, 1866, 1868: oled_data = 16'b1010010010110101;
        1870, 1871, 1872, 1873, 1877, 1878, 1880, 1882, 1883, 1885: oled_data = 16'b1010010010110101;
        1887, 1891, 1892, 1893, 1896, 1898, 1901, 1903, 1957, 1959: oled_data = 16'b1010010010110101;
        1960, 1962, 1964, 1965, 1970, 1971, 1972, 1974, 1975, 1977: oled_data = 16'b1010010010110101;
        1979, 1981, 1982, 1984, 1985, 1990, 1992, 1993, 1995: oled_data = 16'b1010010010110101;
        1614, 1763, 1859: oled_data = 16'b0110101100001111;
        1616: oled_data = 16'b1110111010111011;
        1649, 1940: oled_data = 16'b1110001100001100;
        1650: oled_data = 16'b1111001101001100;
        1655: oled_data = 16'b1111111000111001;
        1656: oled_data = 16'b1111011001111010;
        1658: oled_data = 16'b0110101001001011;
        1660, 1662, 1854, 1856: oled_data = 16'b1110101100001000;
        1661, 1663, 1758: oled_data = 16'b1111001011001000;
        1664, 2044: oled_data = 16'b1100001011001000;
        1665: oled_data = 16'b1010001010001001;
        1666: oled_data = 16'b0101101011001110;
        1667, 1998: oled_data = 16'b1000001110010001;
        1669, 1677, 1683, 1687, 1693, 1696, 1699, 1702, 1705, 1781: oled_data = 16'b1010010001010101;
        1788, 1806, 1862, 1867, 1875, 1881, 1888, 1890, 1895, 1899: oled_data = 16'b1010010001010101;
        1956, 1967, 1969, 1980, 1987, 1989, 1996: oled_data = 16'b1010010001010101;
        1672, 1690, 1708, 1770, 1775, 1777, 1797, 1864, 1869, 1879: oled_data = 16'b1010010001010100;
        1886, 1897, 1961, 1973, 1978: oled_data = 16'b1010010001010100;
        1710, 1809, 1905, 1955: oled_data = 16'b1000110000010010;
        1711, 1954: oled_data = 16'b1000001110010000;
        1712: oled_data = 16'b0111101101001111;
        1713: oled_data = 16'b1011010100110101;
        1742: oled_data = 16'b0101001001001010;
        1743: oled_data = 16'b1000001001001011;
        1744, 1841: oled_data = 16'b1100101011001010;
        1746: oled_data = 16'b1110101100001011;
        1747, 1844, 1941: oled_data = 16'b1111001110001101;
        1750: oled_data = 16'b1111110000010000;
        1751: oled_data = 16'b1111111000111000;
        1752: oled_data = 16'b1111010111111000;
        1753: oled_data = 16'b1110001101001101;
        
        1754, 1937, 2034: oled_data = 16'b0111001001001010;
        1761, 1857: oled_data = 16'b1110001011001000;
        1843: oled_data = 16'b1110001011001010;
        1845: oled_data = 16'b1111110010110010;
        1847: oled_data = 16'b1111110010110001;
        1848: oled_data = 16'b1100001100001100;
        1850: oled_data = 16'b1011001010001001;
        1852, 1950: oled_data = 16'b1111001100001000;
        1858: oled_data = 16'b0011000111001001;
        1935: oled_data = 16'b1101010111111001;
        1936, 2231, 2235, 2237, 2238, 2240, 2242, 2244, 2246, 2248: oled_data = 16'b1011010011110100;
        2250, 2252, 2254, 2256, 2258, 2260, 2262, 2264, 2266, 2268: oled_data = 16'b1011010011110100;
        2270, 2272, 2274, 2276, 2278, 2280, 2282, 2284: oled_data = 16'b1011010011110100;
        1938: oled_data = 16'b1010001010001011;
        1942: oled_data = 16'b1111110011110011;
        1943: oled_data = 16'b1001001100001101;
        1944: oled_data = 16'b1000001010001010;
        1945: oled_data = 16'b1010101010001001;
        1946: oled_data = 16'b1101101011001000;
        1952: oled_data = 16'b1001101001001001;
        1953: oled_data = 16'b0110001001001001;
        1999: oled_data = 16'b0110001011001101;
        2000: oled_data = 16'b1010110010110100;
        2001: oled_data = 16'b1100110111111000;
        2033: oled_data = 16'b0101001001001011;
        2035: oled_data = 16'b1011101010001011;
        2036: oled_data = 16'b1101001011001010;
        2037: oled_data = 16'b1101001100001011;
        2038: oled_data = 16'b1100101101001101;
        2041: oled_data = 16'b1011101010001000;
        2042, 2045, 2047: oled_data = 16'b1100001011001001;
        2043, 2046: oled_data = 16'b1100001010001000;
        2048: oled_data = 16'b0110101000001001;
        2050, 2054, 2057, 2062, 2069, 2072, 2079, 2082, 2086, 2089: oled_data = 16'b1000101111010010;
        2092: oled_data = 16'b1000101111010010;
        2094: oled_data = 16'b0110101011001110;
        2096, 4159, 4570: oled_data = 16'b1110111010111100;
        2132: oled_data = 16'b1100001010001011;
        2190: oled_data = 16'b1001010001010011;
        2226: oled_data = 16'b1101111000111001;
        2227, 2230, 2232, 2234, 2236, 2239, 2241, 2243, 2245, 2247: oled_data = 16'b1010110011110100;
        2249, 2251, 2253, 2255, 2257, 2259, 2261, 2263, 2265, 2267: oled_data = 16'b1010110011110100;
        2269, 2271, 2273, 2275, 2277, 2279, 2281, 2283, 2285: oled_data = 16'b1010110011110100;
        2229: oled_data = 16'b0111101011001100;
        2233: oled_data = 16'b1011010010110100;
        2286: oled_data = 16'b1101010111111000;
        2324: oled_data = 16'b0111001100001101;
        2325: oled_data = 16'b1000101110010001;
        2802, 3106, 3202: oled_data = 16'b1111010111111101;
        2803, 2850, 4174: oled_data = 16'b1011110000011000;
        2804, 2806, 2814, 2822, 2837, 2843, 2852, 4143, 4144, 4146: oled_data = 16'b1011010000011000;
        4150, 4152, 4183, 4191: oled_data = 16'b1011010000011000;
        2805, 2807, 2813, 2821, 2849, 2851, 2853, 4142, 4145, 4151: oled_data = 16'b1011010000010111;
        4158, 4175: oled_data = 16'b1011010000010111;
        2808: oled_data = 16'b1100010011111000;
        2812, 2820, 4149: oled_data = 16'b1110010011111011;
        2815, 4352: oled_data = 16'b1101010111111010;
        2823, 2854: oled_data = 16'b1101010110111010;
        2832, 4141, 4200: oled_data = 16'b1101110011111011;
        2833, 2844, 4184: oled_data = 16'b1011010001010111;
        2836: oled_data = 16'b1110110110111101;
        2838, 2858, 3530, 4147, 4198: oled_data = 16'b1110011001111011;
        2841, 4173: oled_data = 16'b1111011000111101;
        2842, 4190: oled_data = 16'b1100010000011000;
        2848, 4196: oled_data = 16'b1110110100111100;
        2856, 4567: oled_data = 16'b1110110110111100;
        2857: oled_data = 16'b1011110000010111;
        2898: oled_data = 16'b1111110000011110;
        2899, 4575: oled_data = 16'b0101000011001111;
        2900, 2901, 2903, 2909, 2910, 2917, 2918, 2929, 2939, 2945: oled_data = 16'b0011100011001110;
        2947, 2948, 2949, 3049, 3125, 3129, 3139, 3145, 3217, 3221: oled_data = 16'b0011100011001110;
        3235, 3241, 3313, 3317, 3321, 3331, 3413, 3417, 3505, 3509: oled_data = 16'b0011100011001110;
        
        3523, 3582, 3589, 3590, 3611, 3612, 3619, 3625, 4238, 4239: oled_data = 16'b0011100011001110;
        4242, 4246, 4247, 4248, 4254, 4271, 4279, 4280, 4287, 4293: oled_data = 16'b0011100011001110;
        4342, 4389, 4393, 4432, 4438, 4461, 4465, 4469, 4477, 4485: oled_data = 16'b0011100011001110;
        4489, 4534, 4557, 4561, 4565, 4577, 4624, 4641, 4653, 4657: oled_data = 16'b0011100011001110;
        4664, 4665, 4669, 4677, 4681, 4685, 4686, 4720, 4726, 4737: oled_data = 16'b0011100011001110;
        4753, 4757, 4773, 4816, 4822, 4833, 4845, 4849, 4861, 4869: oled_data = 16'b0011100011001110;
        4873, 4912, 4918, 4922, 4941, 4945, 4951, 4952, 4965: oled_data = 16'b0011100011001110;
        2902, 2933, 3043, 3121, 3133, 3225, 3229, 3325, 3421, 4240: oled_data = 16'b0100000011001110;
        4249, 4297, 4442, 4450, 4481, 4630, 4661, 4769, 4826, 4957: oled_data = 16'b0100000011001110;
        4961: oled_data = 16'b0100000011001110;
        2904, 4588: oled_data = 16'b0011001000010001;
        2905, 3715, 5041: oled_data = 16'b1010111101111101;
        2908: oled_data = 16'b1011100101011001;
        2911: oled_data = 16'b0100010000010101;
        2916: oled_data = 16'b1011101001011001;
        2919: oled_data = 16'b0011010001010110;
        2928, 3216, 3408, 4237, 4460, 4488, 4584, 4640, 4652, 4832: oled_data = 16'b1011000111011000;
        4968: oled_data = 16'b1011000111011000;
        2930, 2941: oled_data = 16'b1000011100111101;
        2932, 3412, 3508, 4464, 4752, 4944: oled_data = 16'b1110001111011100;
        2934: oled_data = 16'b0100010101111001;
        2937, 4269, 4277, 4864: oled_data = 16'b1111110010111101;
        2938, 4278, 4286: oled_data = 16'b0101100011010001;
        2940, 2946, 2953, 3025, 3029, 3112, 3337, 3409, 3427, 3581: oled_data = 16'b0011100100001110;
        3601, 3605, 4241, 4288, 4336, 4528, 4585, 4673, 4749, 4761: oled_data = 16'b0011100100001110;
        4765, 4929, 4969: oled_data = 16'b0011100100001110;
        2944, 4484, 4580, 4868: oled_data = 16'b1101101010011100;
        2950, 3513: oled_data = 16'b0011101111010101;
        2952, 3048, 3240, 3336, 3624: oled_data = 16'b1101101101011011;
        2954: oled_data = 16'b0101010110111010;
        2995: oled_data = 16'b1011011010111100;
        2996: oled_data = 16'b0111011001111101;
        2997: oled_data = 16'b0100100111010010;
        2998, 3094, 3286, 3382: oled_data = 16'b0010101100010011;
        2999: oled_data = 16'b0101111100111101;
        3000, 3006, 3013, 3014, 3035, 3045, 4338, 4344, 4367, 4375: oled_data = 16'b0110111100111101;
        4383: oled_data = 16'b0110111100111101;
        3001, 3017, 3095, 3191, 3383, 3575, 5049: oled_data = 16'b1100011100111101;
        3002, 3098, 3290: oled_data = 16'b1111110100111110;
        3003: oled_data = 16'b0111000011010010;
        3004: oled_data = 16'b0101101100010100;
        3005, 3046, 4586, 4778: oled_data = 16'b0111011100111101;
        3007: oled_data = 16'b0101101011010111;
        3008: oled_data = 16'b0100100110010000;
        3009, 3205, 5072: oled_data = 16'b1101011100111101;
        3010, 3298, 3394, 3482: oled_data = 16'b1111110111111101;
        3011: oled_data = 16'b0111000011010011;
        3012: oled_data = 16'b0101101011010100;
        3015: oled_data = 16'b0101001101010110;
        3016, 4377: oled_data = 16'b0100100101010000;
        3024, 3120, 3504, 4296, 4556, 4776, 4844, 4872, 4928: oled_data = 16'b1010100111011000;
        3026, 3602, 4970: oled_data = 16'b0111011100111110;
        3028, 3604: oled_data = 16'b1110001110011100;
        3030, 3222, 3510, 3606, 4946: oled_data = 16'b0011110101111001;
        3032, 4245, 4372, 4756: oled_data = 16'b1100100111011010;
        3033, 4365, 4373, 4381: oled_data = 16'b0100100100001111;
        3034, 4374: oled_data = 16'b0110110111111011;
        3036: oled_data = 16'b0111010110111101;
        3037, 4346, 4558: oled_data = 16'b0100000101010000;
        3038, 4386, 4395: oled_data = 16'b0111010010110111;
        3040: oled_data = 16'b1111011010111100;
        3041: oled_data = 16'b1000111011111101;
        3042, 4376: oled_data = 16'b0110110110111101;
        3044: oled_data = 16'b0011010010110111;
        3050, 3146, 3242, 3338, 4390, 4486, 4582, 4678, 4774, 4870: oled_data = 16'b0100010111111010;
        4966: oled_data = 16'b0100010111111010;
        
        3092: oled_data = 16'b1111110101111110;
        3093, 3189, 3291: oled_data = 16'b0110100010010010;
        3099, 3299: oled_data = 16'b0110000010010010;
        3100, 3190, 3300, 3396: oled_data = 16'b0010101101010100;
        3101, 4542: oled_data = 16'b1110111011111101;
        3103, 3295: oled_data = 16'b1001100010010111;
        3104, 3392: oled_data = 16'b0011100100001111;
        3105, 4261, 5054, 5061: oled_data = 16'b1010011101111101;
        3107, 3203, 3285, 3387, 3477: oled_data = 16'b0110100011010010;
        3108, 3196, 3574: oled_data = 16'b0010101101010011;
        3109, 3301, 3397, 3479: oled_data = 16'b1100111100111101;
        3111: oled_data = 16'b1010000110010111;
        3113, 3209, 3305, 3401, 3677, 3697, 3707, 4339, 5025, 5037: oled_data = 16'b1000011101111110;
        5058, 5065: oled_data = 16'b1000011101111110;
        3122, 3410, 4462, 4834: oled_data = 16'b0111011101111101;
        3124: oled_data = 16'b1110101110011100;
        3126, 3318, 3414, 4466, 4562, 4658, 4754, 4850: oled_data = 16'b0011110110111001;
        3128, 3224, 3320, 4341, 4437, 4468, 4533, 4564, 4629, 4660: oled_data = 16'b1100000111011010;
        4725, 4821, 4917: oled_data = 16'b1100000111011010;
        3130, 4766, 4862: oled_data = 16'b0101111010111100;
        3132, 3138, 3234, 3324, 3330, 3420, 3618: oled_data = 16'b1111101110011110;
        3134, 3422, 4482, 4578, 4674, 4866: oled_data = 16'b0010010010110111;
        3140, 3236, 3332: oled_data = 16'b0100010011110111;
        3144: oled_data = 16'b1101101110011011;
        3188, 4285: oled_data = 16'b1111010101111101;
        3194: oled_data = 16'b1111110011111101;
        3195, 3395: oled_data = 16'b0110000011010010;
        3199: oled_data = 16'b1010000011010111;
        3200, 3400: oled_data = 16'b0011100101001110;
        3201, 3297, 3489, 5009: oled_data = 16'b1010011101111110;
        3204, 3292, 3388: oled_data = 16'b0010001101010100;
        3207: oled_data = 16'b1010000101010111;
        3208, 3296, 3304: oled_data = 16'b0011100101001111;
        3218, 4385, 4394, 4535: oled_data = 16'b0100000101001111;
        3219, 4560, 4576: oled_data = 16'b0101000011010000;
        3220: oled_data = 16'b0100100100010000;
        3226, 3418, 4478, 4958: oled_data = 16'b0101111010111011;
        3228, 4825: oled_data = 16'b1111001110011110;
        3230, 4962: oled_data = 16'b0010010011110111;
        3284, 3476: oled_data = 16'b1111110100111101;
        3287: oled_data = 16'b1100111100111110;
        3303: oled_data = 16'b1010000101010110;
        3312, 4392, 4680: oled_data = 16'b1010100111010111;
        3314, 3315, 3496, 4632, 4655, 4671: oled_data = 16'b0010010000010110;
        3316, 4656: oled_data = 16'b0010001111010101;
        3322: oled_data = 16'b0101111001111100;
        3326: oled_data = 16'b0010010011111000;
        3380, 3572, 4472: oled_data = 16'b1111110101111101;
        3381, 3573: oled_data = 16'b0110100010010011;
        3386: oled_data = 16'b1111010100111101;
        3391: oled_data = 16'b1010000010010110;
        3393, 4273, 5008: oled_data = 16'b1001111101111101;
        3399: oled_data = 16'b1001100101010111;
        3411, 3579, 4532, 4626, 4628, 4637, 4639, 4723, 4728, 4733: oled_data = 16'b1110111100111101;
        4751, 4767, 4954: oled_data = 16'b1110111100111101;
        3416: oled_data = 16'b1100100111011001;
        3426: oled_data = 16'b1111001101011110;
        3428, 3620: oled_data = 16'b0100110011110111;
        3432: oled_data = 16'b1111011001111101;
        3433: oled_data = 16'b1000111001111100;
        3434, 3506, 4334, 4846: oled_data = 16'b0111111100111101;
        3478: oled_data = 16'b0010101100010100;
        3483: oled_data = 16'b0111101101010111;
        3484: oled_data = 16'b0001110001010110;
        3485: oled_data = 16'b1010001111010110;
        3486, 3494, 3515, 4855: oled_data = 16'b1010101111010111;
        3487: oled_data = 16'b1001001001010110;
        3488, 4633: oled_data = 16'b0001110000010110;
        3490, 4189: oled_data = 16'b1111111001111101;
        3491: oled_data = 16'b1000001101010111;
        3492, 4490, 4672: oled_data = 16'b0010010001010110;
        3493: oled_data = 16'b1000110000010111;
        3495: oled_data = 16'b1001101001010110;
        3497, 5014: oled_data = 16'b1000111101111110;
        3512: oled_data = 16'b1101101111011011;
        3514: oled_data = 16'b0100110001010111;
        
        3516, 4856: oled_data = 16'b1010001010010111;
        3517: oled_data = 16'b0101101110010101;
        3518: oled_data = 16'b0001111000111011;
        3522: oled_data = 16'b1111101110011101;
        3524: oled_data = 16'b0100010011111000;
        3528: oled_data = 16'b1110110101111100;
        3529: oled_data = 16'b1010110000010110;
        3580: oled_data = 16'b1011000110011001;
        3583: oled_data = 16'b0011110000010110;
        3584, 3614, 3671, 4453, 5070: oled_data = 16'b1110011100111101;
        3588: oled_data = 16'b1010101010011001;
        3591: oled_data = 16'b0010110001010110;
        3592, 3669: oled_data = 16'b1101111100111101;
        3600, 4748, 4940: oled_data = 16'b1011000111010111;
        3609, 4949: oled_data = 16'b1110110011111110;
        3610: oled_data = 16'b0101000011010001;
        3613, 4874: oled_data = 16'b0111111101111101;
        3626: oled_data = 16'b0100110111111010;
        3670, 3678, 3687, 4738, 4930, 5048, 5071: oled_data = 16'b0111111101111110;
        3679: oled_data = 16'b1000111101111101;
        3685, 3722, 4953: oled_data = 16'b1001011101111101;
        3686, 3708: oled_data = 16'b0111111110111110;
        3698, 4304: oled_data = 16'b1011111101111101;
        3701: oled_data = 16'b1010111100111101;
        3702, 3716, 4357, 5019, 5042, 5053: oled_data = 16'b1001011101111110;
        3706: oled_data = 16'b1100111101111101;
        3709, 5038, 5046, 5057, 5066: oled_data = 16'b1011111100111101;
        3721, 5018: oled_data = 16'b1010111101111110;
        4153: oled_data = 16'b1011010010111000;
        4155, 4440: oled_data = 16'b1111111100111110;
        4157: oled_data = 16'b1110010101111100;
        4163: oled_data = 16'b1101010001011010;
        4164, 4176: oled_data = 16'b1011110010111000;
        4181, 4353: oled_data = 16'b1111111000111101;
        4182: oled_data = 16'b1100010000011001;
        4192, 4197, 4201: oled_data = 16'b1011010001011000;
        4206: oled_data = 16'b1100110000011001;
        4207: oled_data = 16'b1100010100111001;
        4243: oled_data = 16'b0100110101111001;
        4250, 5062: oled_data = 16'b1001111101111110;
        4251, 4340: oled_data = 16'b1111111101111101;
        4252, 4445: oled_data = 16'b1111111101111110;
        4253, 4668: oled_data = 16'b1100001010011010;
        4255: oled_data = 16'b0110111010111011;
        4259: oled_data = 16'b1001000100010110;
        4260: oled_data = 16'b0011100111010000;
        4270, 4865: oled_data = 16'b0100000011001111;
        4272: oled_data = 16'b0011100110010000;
        4281: oled_data = 16'b1010011100111101;
        4289: oled_data = 16'b1000111100111110;
        4292: oled_data = 16'b1110001010011100;
        4294: oled_data = 16'b0101010111111010;
        4298: oled_data = 16'b1000011101111101;
        4302, 4494, 4878, 4974: oled_data = 16'b0111100010010100;
        4303, 4399, 4687, 4879: oled_data = 16'b0011001010010010;
        4333: oled_data = 16'b1111011001111100;
        4335: oled_data = 16'b0110010001011001;
        4337, 4474: oled_data = 16'b0011011000111011;
        4343: oled_data = 16'b0100011001111011;
        4345, 4384: oled_data = 16'b0110110111111101;
        4347: oled_data = 16'b1000010010110111;
        4348, 4434: oled_data = 16'b1111011101111110;
        4349: oled_data = 16'b1101001111011011;
        4350: oled_data = 16'b0011101011010011;
        4351: oled_data = 16'b0101010011111001;
        4354: oled_data = 16'b1100010001011001;
        4355: oled_data = 16'b1001000111010110;
        4356, 4670: oled_data = 16'b0010001110010100;
        4364: oled_data = 16'b1011001000011000;
        4366: oled_data = 16'b0111011010111101;
        4368: oled_data = 16'b0110110101111100;
        4369: oled_data = 16'b0100000100001111;
        4370: oled_data = 16'b1000010101111001;
        4378: oled_data = 16'b0111110010110111;
        4380, 4956: oled_data = 16'b1100001011011010;
        4382: oled_data = 16'b0111010111111011;
        4388, 4772, 4964: oled_data = 16'b1101101010011011;
        4398, 4590: oled_data = 16'b0111100010010011;
        4400, 4592: oled_data = 16'b1011011100111110;
        4431, 4527, 4623, 4719, 4815, 4911: oled_data = 16'b1100101011011010;
        4433, 4721: oled_data = 16'b0101011001111011;
        4439, 4758: oled_data = 16'b0111111010111011;
        4441, 4921: oled_data = 16'b1111101111011110;
        4443, 4731, 4762, 4923: oled_data = 16'b0100010010110111;
        
        4444: oled_data = 16'b1111011101111101;
        4446: oled_data = 16'b1100111000111110;
        4447, 4536, 4537: oled_data = 16'b0101000100010000;
        4448: oled_data = 16'b0011101110010101;
        4449: oled_data = 16'b1110010010111110;
        4451, 4827: oled_data = 16'b0011110010110111;
        4452: oled_data = 16'b1100011100111110;
        4470: oled_data = 16'b1000011001111011;
        4473: oled_data = 16'b0100110000010110;
        4476, 4572, 4764, 4860: oled_data = 16'b1100001010011001;
        4480: oled_data = 16'b1111110010111110;
        4491: oled_data = 16'b0010010001010111;
        4492: oled_data = 16'b1010010001010110;
        4493: oled_data = 16'b1111111010111101;
        4495, 4591, 4783, 4975: oled_data = 16'b0010101010010010;
        4496, 4688, 4880, 5015: oled_data = 16'b1011011101111101;
        4529, 4913: oled_data = 16'b0101111001111011;
        4538: oled_data = 16'b0110111010111100;
        4539, 4642, 4682, 4750, 4942: oled_data = 16'b0111011101111110;
        4543: oled_data = 16'b1010110111111100;
        4544: oled_data = 16'b0100101111010111;
        4545: oled_data = 16'b0101000101010000;
        4546: oled_data = 16'b0111011000111100;
        4547: oled_data = 16'b0110011100111101;
        4559: oled_data = 16'b0101000100001111;
        4566, 4662, 4823, 4919: oled_data = 16'b0111111001111011;
        4568: oled_data = 16'b1101010100111011;
        4569: oled_data = 16'b1101110100111010;
        4573, 4730, 4777: oled_data = 16'b0100000100001110;
        4574: oled_data = 16'b0011100101010000;
        4581: oled_data = 16'b0100000011001101;
        4587: oled_data = 16'b1001100101010110;
        4589: oled_data = 16'b1000111010111101;
        4625: oled_data = 16'b0101011001111100;
        4631: oled_data = 16'b0010001110010101;
        4634: oled_data = 16'b0110110001010111;
        4635: oled_data = 16'b1100110110111010;
        4654: oled_data = 16'b0010010000010101;
        4663: oled_data = 16'b1011000100011000;
        4666: oled_data = 16'b0101110010110111;
        4676: oled_data = 16'b1101101001011100;
        4684: oled_data = 16'b1000010101111101;
        4727: oled_data = 16'b0111011001111011;
        4729: oled_data = 16'b1110101111011110;
        4736: oled_data = 16'b1010101000011000;
        4759: oled_data = 16'b1110010100111100;
        4760: oled_data = 16'b0100110101111011;
        4768, 4960: oled_data = 16'b1111010010111110;
        4770: oled_data = 16'b0010010010111000;
        4780: oled_data = 16'b1111010110111101;
        4781: oled_data = 16'b0110110011111000;
        4782: oled_data = 16'b0011101000010001;
        4784, 4976: oled_data = 16'b1011011101111110;
        4817: oled_data = 16'b0101011010111011;
        4848: oled_data = 16'b1110101111011100;
        4852: oled_data = 16'b1101110000011011;
        4853: oled_data = 16'b0010101111010101;
        4854: oled_data = 16'b0101110001010111;
        4857: oled_data = 16'b0100101110010101;
        4858: oled_data = 16'b0011010111111010;
        4877: oled_data = 16'b1111011010111101;
        4950: oled_data = 16'b0101100011010000;
        5026: oled_data = 16'b1011011100111101;
        5047: oled_data = 16'b1000011110111110;
        default: oled_data = 16'b0000000000000000;
        endcase

    end endmodule
